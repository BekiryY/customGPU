//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.03 (64-bit)
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Wed Dec 10 21:11:32 2025

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [15:0] ad;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire [30:0] prom_inst_2_dout_w;
wire [0:0] prom_inst_2_dout;
wire [30:0] prom_inst_3_dout_w;
wire [0:0] prom_inst_3_dout;
wire [30:0] prom_inst_4_dout_w;
wire [1:1] prom_inst_4_dout;
wire [30:0] prom_inst_5_dout_w;
wire [1:1] prom_inst_5_dout;
wire [30:0] prom_inst_6_dout_w;
wire [1:1] prom_inst_6_dout;
wire [30:0] prom_inst_7_dout_w;
wire [1:1] prom_inst_7_dout;
wire [30:0] prom_inst_8_dout_w;
wire [2:2] prom_inst_8_dout;
wire [30:0] prom_inst_9_dout_w;
wire [2:2] prom_inst_9_dout;
wire [30:0] prom_inst_10_dout_w;
wire [2:2] prom_inst_10_dout;
wire [30:0] prom_inst_11_dout_w;
wire [2:2] prom_inst_11_dout;
wire [30:0] prom_inst_12_dout_w;
wire [3:3] prom_inst_12_dout;
wire [30:0] prom_inst_13_dout_w;
wire [3:3] prom_inst_13_dout;
wire [30:0] prom_inst_14_dout_w;
wire [3:3] prom_inst_14_dout;
wire [30:0] prom_inst_15_dout_w;
wire [3:3] prom_inst_15_dout;
wire [30:0] prom_inst_16_dout_w;
wire [4:4] prom_inst_16_dout;
wire [30:0] prom_inst_17_dout_w;
wire [4:4] prom_inst_17_dout;
wire [30:0] prom_inst_18_dout_w;
wire [4:4] prom_inst_18_dout;
wire [30:0] prom_inst_19_dout_w;
wire [4:4] prom_inst_19_dout;
wire [30:0] prom_inst_20_dout_w;
wire [5:5] prom_inst_20_dout;
wire [30:0] prom_inst_21_dout_w;
wire [5:5] prom_inst_21_dout;
wire [30:0] prom_inst_22_dout_w;
wire [5:5] prom_inst_22_dout;
wire [30:0] prom_inst_23_dout_w;
wire [5:5] prom_inst_23_dout;
wire [30:0] prom_inst_24_dout_w;
wire [6:6] prom_inst_24_dout;
wire [30:0] prom_inst_25_dout_w;
wire [6:6] prom_inst_25_dout;
wire [30:0] prom_inst_26_dout_w;
wire [6:6] prom_inst_26_dout;
wire [30:0] prom_inst_27_dout_w;
wire [6:6] prom_inst_27_dout;
wire [30:0] prom_inst_28_dout_w;
wire [7:7] prom_inst_28_dout;
wire [30:0] prom_inst_29_dout_w;
wire [7:7] prom_inst_29_dout;
wire [30:0] prom_inst_30_dout_w;
wire [7:7] prom_inst_30_dout;
wire [30:0] prom_inst_31_dout_w;
wire [7:7] prom_inst_31_dout;
wire dff_q_0;
wire dff_q_1;
wire mux_o_0;
wire mux_o_1;
wire mux_o_3;
wire mux_o_4;
wire mux_o_6;
wire mux_o_7;
wire mux_o_9;
wire mux_o_10;
wire mux_o_12;
wire mux_o_13;
wire mux_o_15;
wire mux_o_16;
wire mux_o_18;
wire mux_o_19;
wire mux_o_21;
wire mux_o_22;

LUT3 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15])
);
defparam lut_inst_0.INIT = 8'h02;
LUT3 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15])
);
defparam lut_inst_1.INIT = 8'h08;
LUT3 lut_inst_2 (
  .F(lut_f_2),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15])
);
defparam lut_inst_2.INIT = 8'h20;
LUT3 lut_inst_3 (
  .F(lut_f_3),
  .I0(ce),
  .I1(ad[14]),
  .I2(ad[15])
);
defparam lut_inst_3.INIT = 8'h80;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hC8F300ACB0B4B4896FF873435E56A804B7FFFF18000064726E8B451A6ADF9AD0;
defparam prom_inst_0.INIT_RAM_01 = 256'hA4DB7FEC7D81831931634F6EAFF1836772AD10093FFFF7100000C1C4DEBE9008;
defparam prom_inst_0.INIT_RAM_02 = 256'hC0031C6CB465D71C3FF8EABB62CD27719FFE7A647251601B7FFFE71FE001831C;
defparam prom_inst_0.INIT_RAM_03 = 256'h7F8063800006738D171A01E3E48E2C1A45A5E2DB40238DBE9FCABFDA7FFFC73F;
defparam prom_inst_0.INIT_RAM_04 = 256'h2F550096FF00E300000C8F5CD16CEBD4DAE35D920B341E8F80389654291A7F92;
defparam prom_inst_0.INIT_RAM_05 = 256'hFE312C0309B601A7FFFEE3FE0018389B55D22863FA70469616D38220FFCFD357;
defparam prom_inst_0.INIT_RAM_06 = 256'h59B28C33FDC34D27936C036FFFFCE3FC00306314BB2FF389B47173A62C484EFD;
defparam prom_inst_0.INIT_RAM_07 = 256'h90CC812E4F5B53586698C472A8E0E69C99847387FF98E62D96BFFEDA38E6A36C;
defparam prom_inst_0.INIT_RAM_08 = 256'h5AF46D3AB9EDE40C9AC8C851CD30CDD551C1CD33618E7F1FFE318C5B2D7EBCB7;
defparam prom_inst_0.INIT_RAM_09 = 256'hC338F16CB5C00921F8F599E506293F871A7CEE2AA3839A6D18E31CFFF8E618B6;
defparam prom_inst_0.INIT_RAM_0A = 256'h47E38E001C63E2D96BAE4B689821BDCDBF2560BCF4CE0395470734E4CC3C73FF;
defparam prom_inst_0.INIT_RAM_0B = 256'h1C1CD3D3711C3000F10CC5B2D7FDDBC8185BA3EBC5259663E9E3F8AA8E0E6996;
defparam prom_inst_0.INIT_RAM_0C = 256'hA61DBAAA3839A66839C7E7FFC6318B65AFC7921C1CC7BFC9F7E1020ED3380A55;
defparam prom_inst_0.INIT_RAM_0D = 256'h571B44E34F1FD55470734CB23CE38FFF1CE316CB5E8DA48A3DAEE2127CF18239;
defparam prom_inst_0.INIT_RAM_0E = 256'hBE2AEDE612D55341C59487E8C73A3A0315EAA739C6392769077FF99D5EFC9CA1;
defparam prom_inst_0.INIT_RAM_0F = 256'h1DE0029A34D0F173896DB341C5C90691CE73BAE1DAC8FE718C7244D20EF00388;
defparam prom_inst_0.INIT_RAM_10 = 256'hF1F2C6883BC01095275468C0C3449961D477A811FCE6D15CB8FCFCE198F543C4;
defparam prom_inst_0.INIT_RAM_11 = 256'h58FFF3F1E3EAD19077FF9416715E2E37A79565B1D35BC0B9F9F3078CB4E5B9F1;
defparam prom_inst_0.INIT_RAM_12 = 256'hE7A797F4A51AE730C774E520EFFF72AA8D6A6DA4E4C592798D25DFB8F3B5F201;
defparam prom_inst_0.INIT_RAM_13 = 256'h9B20D239CE773F3BA7EBCE318E5C9A41DE00A3B7E73FF949FE2EC938A390FD18;
defparam prom_inst_0.INIT_RAM_14 = 256'h79D34C3396D1023B9DA2F7CC5CD39C731CA97483BC005B6EB9F03447C5A22C38;
defparam prom_inst_0.INIT_RAM_15 = 256'hB6BA407F8638C205627A0A1FFBDA152FB4E0AC8C9D551DFC41279A9C691E9620;
defparam prom_inst_0.INIT_RAM_16 = 256'hA49203A0C0FB152948E38D7666A4233F01F02A2897C439A9624B2BF822405B86;
defparam prom_inst_0.INIT_RAM_17 = 256'h1568D0420903183CCB5B7245E39E23A26437E534F8D7CBF13384BB269B6B880E;
defparam prom_inst_0.INIT_RAM_18 = 256'hBEE3F165972C5EF9923210C0E3BC7F1F4E39C08021505E2D752F6425B8C7494B;
defparam prom_inst_0.INIT_RAM_19 = 256'h69423C919C6CB0D38BE7B64C24799CDBC74E889E71C7089B795F789592B4F834;
defparam prom_inst_0.INIT_RAM_1A = 256'h7205DA161C05E122FBC8CD2CE8757F64485B0EAFA54D1AA5C718E335DE69A97E;
defparam prom_inst_0.INIT_RAM_1B = 256'h71C62A0322FAE99B5A5B59BE0CB700DB45629BCC90F4679E1F206A391C710284;
defparam prom_inst_0.INIT_RAM_1C = 256'h297143E63822EE258B1455EE5B6128D1BCB06E5AA9326A20F1CA738852B6040C;
defparam prom_inst_0.INIT_RAM_1D = 256'hD38A0B9083BA436C7818B84B05A189C6D423C1A9499FDE9552E4D441E19B981F;
defparam prom_inst_0.INIT_RAM_1E = 256'h76535107B1AC000F0553E158EB11B4840521EB6E6792C3558BE7CD8AB549A883;
defparam prom_inst_0.INIT_RAM_1F = 256'h75934BAAAAA6A20F31DDDCD71849E0F1D4950E92B1E47540DC2F4680A8DC4D15;
defparam prom_inst_0.INIT_RAM_20 = 256'h3F6F1AA70792DB55064D441E397504DB9E87AB63A554ADEFC7B8E38E7D5C8D37;
defparam prom_inst_0.INIT_RAM_21 = 256'h903F1218587834898725D2AA5C9A883D316D321E883383C71A2D47B76BA0D51D;
defparam prom_inst_0.INIT_RAM_22 = 256'h813A908208C063414FA06B0FBB35A156B935107A72B4690C09DDD98F03AB0860;
defparam prom_inst_0.INIT_RAM_23 = 256'h81C4CE01C9C2AC8FF58C7788DB4DA2A07F4C5D5E9D97794320BD197A2FEA0B1C;
defparam prom_inst_0.INIT_RAM_24 = 256'h855EF910C11A90303BA559EE6A469998976C803E7E962ABD3B2EF246431C29F1;
defparam prom_inst_0.INIT_RAM_25 = 256'hECBBF5D909EC6AE186375D9F4F4AB0F5E0DE09D026903129DD3CB57A765DE6CC;
defparam prom_inst_0.INIT_RAM_26 = 256'h74F2D5E9D977E4B277F4CEC241B7729613D56D20278ACB8BCB71D26CBA7E6AF4;
defparam prom_inst_0.INIT_RAM_27 = 256'hA24DF3B7E95DABD3B2EF286467DAF6517119DF9B0E2A97D42E471CD6C2D5C3BD;
defparam prom_inst_0.INIT_RAM_28 = 256'h7F559BEA7B02774FD27557A765DE68C9AA4155A44DF9D1A51B551AF7D055F166;
defparam prom_inst_0.INIT_RAM_29 = 256'h3D546E79FDA66D18D1C7E57FA5C6AF4ECBBCD991EE279CD9012EAC6FFCAA0C4E;
defparam prom_inst_0.INIT_RAM_2A = 256'hC18FC3F7ED5765855B4C7197D351FE71D05822690BA9C4F67D7B827FE14DD7E7;
defparam prom_inst_0.INIT_RAM_2B = 256'h7B2BFAD0ED26CF3AEAA292CAACBCC1BBE4DD43EB2BB8AC52136389EC738E07A1;
defparam prom_inst_0.INIT_RAM_2C = 256'h5D4E278C21EDB71E2D73E6CF3557D325D2D8075AD0DF09F4768AF464314713DC;
defparam prom_inst_0.INIT_RAM_2D = 256'hB8C52C10C51C4F0E557BC631E24694366A960E9D1A1A5B10FB9494F95D082C88;
defparam prom_inst_0.INIT_RAM_2E = 256'hC438691AD8924D216D389E8F349D080E44AE56715518FDE8CBB4E5F460CD38A6;
defparam prom_inst_0.INIT_RAM_2F = 256'hB798ED8406DAF965C741CA4264713D8EB2F859706B3DA006AA18AB8B2CFC33FC;
defparam prom_inst_0.INIT_RAM_30 = 256'hAA8220AA4E3B6D76CFE902CACA1A9C8608E27B8F2CE02F1FA4F0804155653155;
defparam prom_inst_0.INIT_RAM_31 = 256'h0DD17346FBA0049384899D5E043C992D220575334F19179FC2481F8CC4F2DFF6;
defparam prom_inst_0.INIT_RAM_32 = 256'h8FFEEAD3B955560F98DFF67366FC8A03F5F401A84D22EB661E33230982CF88DE;
defparam prom_inst_0.INIT_RAM_33 = 256'hB8F778C39484E082F94B42AB2B5FF0008FCB3A5CDD3013483B40D7E8A3968193;
defparam prom_inst_0.INIT_RAM_34 = 256'h5A6CA05F0C258E73C5BB77409AD2C6519E401C9F4B4E5B73B145DD13CF955665;
defparam prom_inst_0.INIT_RAM_35 = 256'hAD200B2EF7AA8668AF22E3F1D0005935439134CF3A7FC6B0493F59071760D5AE;
defparam prom_inst_0.INIT_RAM_36 = 256'hFD40C936041EF83C965D7EC2E66870703F83FA504380F314E6FF72F9557FDE84;
defparam prom_inst_0.INIT_RAM_37 = 256'h9003FDFD33ADDA186B28CEA8709AFD0560D0727014AEAC30D0F3F60977FF9D56;
defparam prom_inst_0.INIT_RAM_38 = 256'h3E763B936491BCB4D550FCF7A3AA76B9D165D7F0E497FC7230946C10B7FF96E5;
defparam prom_inst_0.INIT_RAM_39 = 256'h1913DAA0ADFE30CE93E8197D7EB4435E6707169092CB2FE5892FF8038C4871EF;
defparam prom_inst_0.INIT_RAM_3A = 256'hE4803FEE2FB19C21C0FE217FB5E67B72572A21E61BD066624594FFCE72401007;
defparam prom_inst_0.INIT_RAM_3B = 256'h962C7F46C97FBFDC612971D9998E2A2205E53FCDDB9EBDCEC51649664B317FB8;
defparam prom_inst_0.INIT_RAM_3C = 256'h8592A0B02C78FE1C92FF0038F9C6488BF80672D50ED2AF3E4F5AC225A6A98854;
defparam prom_inst_0.INIT_RAM_3D = 256'h669DA0997EBB95165965FCA125FF00716D0BEB0C16C7081736CC66055A310B20;
defparam prom_inst_0.INIT_RAM_3E = 256'h36B0CE0585A83CF96A423284B2DFF9CA480200E37A7B5F794DC65D662BA364A0;
defparam prom_inst_0.INIT_RAM_3F = 256'hE97AA3B2497D9BF4D4BD3B177DBAE8A7FDD6952E8FFC01C6B1E0E56AC7CCD0C3;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hF2542B7F07E2453120E1511FEF19BC778A0917EFFBAD2FF5D00807FFFD2381A8;
defparam prom_inst_1.INIT_RAM_01 = 256'h7FE01FE013A7053A06B179C4E5AE851F1FB909064E1B073FF75A5FF5C0100FFF;
defparam prom_inst_1.INIT_RAM_02 = 256'hDD69001F003FC00014F7C125A8153FCC769B7F853807795EFEE6BB7FEEB496B4;
defparam prom_inst_1.INIT_RAM_03 = 256'hD1950AFFBAD224C1FF7F807FAE2340CC5D553786972F624D061445EE1DEC69FF;
defparam prom_inst_1.INIT_RAM_04 = 256'hFD4DAFEFDF93D9FF75A5FEBC0100FFFFF7A17DE9F355E5F0379DC5C77DEDEF3D;
defparam prom_inst_1.INIT_RAM_05 = 256'h5E1B33CF9971A88A927143FEEB4BFCF80201FFFE8F5963CB6E5DCA3D849973C2;
defparam prom_inst_1.INIT_RAM_06 = 256'h3CA00E640F8107E4EDC074A93E491FFDD720070EAC03FC00279E3F7476A891CE;
defparam prom_inst_1.INIT_RAM_07 = 256'hDD22A62ED9A2DE193BEAC6D623296C9D273B2FFBAE400C5DBF1E9B4945312FCC;
defparam prom_inst_1.INIT_RAM_08 = 256'h5C7A7B78993CCC35FADA3F842A7C36F75D9D42764939DFF757FFF8C5DE3D3C9B;
defparam prom_inst_1.INIT_RAM_09 = 256'h047F9C5538F4E586227FC2D105E05A7BD3FD55DD2ACB9DF283F97FEE86FFC5B5;
defparam prom_inst_1.INIT_RAM_0A = 256'hE4ACFFBAE400E955F1E99231149B5E93A50CAD13D24658E544556C3D1421FFDD;
defparam prom_inst_1.INIT_RAM_0B = 256'hFACB3B0D4343FF75CC018F17E3D3695933AC76916C9D058BB1D8CDBB2D64E599;
defparam prom_inst_1.INIT_RAM_0C = 256'h043FE848EDE044CC377FFEEBDC031EABC7A7960C9AC48B0B0453228E4E9199F0;
defparam prom_inst_1.INIT_RAM_0D = 256'hC56BAA87099A740ED0C76085AE334AF4A167AA6B8F4F6E76ADF7ED2ADDBEDCF2;
defparam prom_inst_1.INIT_RAM_0E = 256'hE528223187C2497BA19DD5787B9842C10AE6C5E942C2C4D1A63FF830D5420E8B;
defparam prom_inst_1.INIT_RAM_0F = 256'h839FEA5283481E96FCFCFCC70BA8C3F900FBD00A40648BD2859A69A248EFF94B;
defparam prom_inst_1.INIT_RAM_10 = 256'h165626B2CE3FCC177A9A6082011CC11FC43F37E0DDF70FF2CC6597A50B02134D;
defparam prom_inst_1.INIT_RAM_11 = 256'h57695E942CF34D69F1FF8727F4B4B54133371AD6EF94AD109E8F355BC2EDAF4A;
defparam prom_inst_1.INIT_RAM_12 = 256'h62F82BA9A258BD2858189A36C7FF93BB9DFD2DFA505B4C55E6863345B0DF0E0D;
defparam prom_inst_1.INIT_RAM_13 = 256'h77D80AD7DAEDA5A7E0917A50B14D34491DFFC322B17CDCE9E604510A50100C0A;
defparam prom_inst_1.INIT_RAM_14 = 256'h02C1E9E5BB5FBC5829F82FB3EE3EF70360A2A0B073FF1A24B9F6DC421800CA2C;
defparam prom_inst_1.INIT_RAM_15 = 256'h49DE5A6A11A7EA8B90E4EF77E3BB30140C78EA96C1C74B840A6A6E8E41DA33CF;
defparam prom_inst_1.INIT_RAM_16 = 256'hBD928F24AFE19E16765879E4CC3A8B9274C9B0707634E3228D65D18BDD948131;
defparam prom_inst_1.INIT_RAM_17 = 256'hCA69DC64D378EA4A103E3404E9F2CD3C76473BE69BFE50BFCE0847E4FAEAF9E6;
defparam prom_inst_1.INIT_RAM_18 = 256'hC75EE46C1455C77F51F0C35992030F9026E9F9A8329D4EC6BDE4DC4D07287B7D;
defparam prom_inst_1.INIT_RAM_19 = 256'h3147F17DCF1D52D8BA49F3EC136BFDA12AEED0A35CDE1D4ABDDADCB68F2B087F;
defparam prom_inst_1.INIT_RAM_1A = 256'h340B2F93311760B3C63C24917C92315626641215BA5D1812752BDB4D7381C75C;
defparam prom_inst_1.INIT_RAM_1B = 256'h6A2B11D9502898772004020E4B6D4907BF1C3AB2CB886087FB631EAACB61EE30;
defparam prom_inst_1.INIT_RAM_1C = 256'h0ECDC511F28673C7473798AD4653C78C96D2920E6E7EA49D38E534DF6B44D76A;
defparam prom_inst_1.INIT_RAM_1D = 256'hB1ECBE89CD0E687B44DDBE5B21A051A714AE0D5B6DA3640199E262C6A70EC37F;
defparam prom_inst_1.INIT_RAM_1E = 256'h9C0C4B10B8DC81BA9BD8E01A1A8A9FC42908F5F1030E0BAD9B558802071E048E;
defparam prom_inst_1.INIT_RAM_1F = 256'h6DE020F7F3ECF4AA9C70812BA427487FF87C0FC588F75AF9F87D601236F21069;
defparam prom_inst_1.INIT_RAM_20 = 256'hC8A53992DA1241DDCF1DCBE60EC3FF729A54EC98938CEA99F04B315B59BECE29;
defparam prom_inst_1.INIT_RAM_21 = 256'h14BE09C164351B2DB46480B31EFCD201E3DA3A1F7FFEC2A9956DF6900FA71AF8;
defparam prom_inst_1.INIT_RAM_22 = 256'h2F5B663E570C117757A00F4C308B2703A2BA5B031D5AF6DC3E58132986812E4B;
defparam prom_inst_1.INIT_RAM_23 = 256'h79F9AAD74490B978F2ED857164F5BF9BF1128F6247D4A69FFAA23083AA89A2A5;
defparam prom_inst_1.INIT_RAM_24 = 256'hE5C2711869676B80E2F5ECD9B244765571C4C2F7E2317CDAA7CC8CBFF7499DBD;
defparam prom_inst_1.INIT_RAM_25 = 256'h8CCC74C02AFAF6921BDD8B8A0DAB12BE95216FE246B9E3900466DF4919A0E59F;
defparam prom_inst_1.INIT_RAM_26 = 256'h1174DB24EC92360069E34A0A0FC7710918462A0D598107A5CAE3B2DF88AAA56D;
defparam prom_inst_1.INIT_RAM_27 = 256'h778C937E2251A45CED4797FF5551CE8D491BF13041CE942574B699760357DE40;
defparam prom_inst_1.INIT_RAM_28 = 256'h16BCA2888F9D2AF446ABBEAD290393FE49F868E8C337BFF4CAB253CA293574C6;
defparam prom_inst_1.INIT_RAM_29 = 256'h42FB295D3DD103C5588BA6891476B37EB545B3FC9326D5BEA615F8502DAF64CD;
defparam prom_inst_1.INIT_RAM_2A = 256'h6F89E0D07A98453641F9ED538FF8B7B228EC891DB08410C79A5B74C9A4E95BFA;
defparam prom_inst_1.INIT_RAM_2B = 256'h7BF0B316AEA5BA2EC6B9B1BE63B408D2C26E8CE451DF0CD69AAFD0EF322C47A9;
defparam prom_inst_1.INIT_RAM_2C = 256'hB0C0863CEB921EC95C0CA025291AEA88EEC3C55155E07788A3A325BE9A92DC7E;
defparam prom_inst_1.INIT_RAM_2D = 256'h8E99916EE00173F982B3FF9213ADDBB06FEE6EE4484B342DEDF5BF914755488B;
defparam prom_inst_1.INIT_RAM_2E = 256'h63B5D0451D9513C4454238F361A904A4B9EFE68D4E312E0DFE90E5D32EF42422;
defparam prom_inst_1.INIT_RAM_2F = 256'h96FB97D90C17608A3BD5BB1946FB1FE76471C9EE9006748DAD1F2FDAB7B4BBEC;
defparam prom_inst_1.INIT_RAM_30 = 256'h60B9703D979E89282315BB9200EA6C48EC0B9FCF01D07104D62F65EA7B58191F;
defparam prom_inst_1.INIT_RAM_31 = 256'hB01A4CE93E828314DEB2B46EA3D2521792C1AE4FDB6C99B2B5265FBC3C18D9CB;
defparam prom_inst_1.INIT_RAM_32 = 256'h6379807BAE03F98483732DE0079A76E3DF85E537DC4340359F4DB96B329351DC;
defparam prom_inst_1.INIT_RAM_33 = 256'h8FA5F2C9E1CE81282706F38905D194DDE2E70B73A1D9235007534596A7459A64;
defparam prom_inst_1.INIT_RAM_34 = 256'h154DD4069D341678601578CE450DB1020B864350FD2556E1B56E6B5FF5268549;
defparam prom_inst_1.INIT_RAM_35 = 256'hC380437A55653462EE96340F38D456EE617A739317A376C7F8EE45C04E8A7240;
defparam prom_inst_1.INIT_RAM_36 = 256'h8E7D55037558A6FFAB17801983972D8587E2908B6FC88527D1AFCA088A619478;
defparam prom_inst_1.INIT_RAM_37 = 256'hDFC60C42886699B35BCB8A14552E4E2CE1A64EB46BAE9A4E316AF4905E6D3019;
defparam prom_inst_1.INIT_RAM_38 = 256'h7C9CCC50F7BAD5420D4B3DF7888FD4213878062E80174D3878C200CAB1262AE2;
defparam prom_inst_1.INIT_RAM_39 = 256'h055E6A0D061987540C7AF2407222795A25BD685071D0036790268E5236DB825E;
defparam prom_inst_1.INIT_RAM_3A = 256'hBF45962DB461E5948AE228D6EAC79BC88226A823D3BFD0B416A002E113C489B3;
defparam prom_inst_1.INIT_RAM_3B = 256'hA1FF8F7532E9D95FBFEF3EE7DCD1A6D29D0B4E88E7E588454D52215BB8FFFA8B;
defparam prom_inst_1.INIT_RAM_3C = 256'h0C6485F91DFF334102C9A32D75AB4447777B1A5AE51A9757C54770987B5542E5;
defparam prom_inst_1.INIT_RAM_3D = 256'h95708E9E406908FA3A01B53524D18A5B5FE8C4CFEF99CA0BDDA0B39AA5C7E094;
defparam prom_inst_1.INIT_RAM_3E = 256'h5FBA5346AFEDEC8D2363C6DEBC0117DA68B1347FA57DC1456056CA97A25C1A2B;
defparam prom_inst_1.INIT_RAM_3F = 256'hF91FD6E5764B19E5B14A122CA6C5AA53C7F800180679758D52143A651F6813B6;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[30:0],prom_inst_2_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 1;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hF00132572FC82D3BE45318767F5779886D91D02AEFF005731C72ACA90D69988A;
defparam prom_inst_2.INIT_RAM_01 = 256'h8C34FBE4E41CDAEAD31F627EB9EA04704688064F9B21D8B5FFE00E839C7568DB;
defparam prom_inst_2.INIT_RAM_02 = 256'h00003BA50E2A4F0B41B962C0E5DFCB083D757AE5CA068DD8B670B163C0001B71;
defparam prom_inst_2.INIT_RAM_03 = 256'hD8B54A50FF0004D88F24778861D2B6E7E0BE7646FB58287267847E596C7181E3;
defparam prom_inst_2.INIT_RAM_04 = 256'h2B908AF9B07B6F0DFE00D7438F5584DC99A93BB9C37ADD41F6FA8DE0D8407484;
defparam prom_inst_2.INIT_RAM_05 = 256'h549A4B17F6A6B5A5F0142923FC00A7538EAA99D4FD7423BFB909B58D2EBE5E1A;
defparam prom_inst_2.INIT_RAM_06 = 256'h07D7656B88B94E876265A15A7820055F19C60FE9249AC6CC0A57EE40810C4DDB;
defparam prom_inst_2.INIT_RAM_07 = 256'h778ED48F0412D56711CE932D14D2159B57C1954181CCD1524961633A949E7A1B;
defparam prom_inst_2.INIT_RAM_08 = 256'h0B10AD5950A1C22A8DFD8FA98146AA6BAEECCC617F5836E1D8F5312486917F59;
defparam prom_inst_2.INIT_RAM_09 = 256'hE3FFE31265EDB30F22C77AE805B7BF4977F2D070A78E1803A0FC2A460E26EDC9;
defparam prom_inst_2.INIT_RAM_0A = 256'h0485AB8E30C89A24D39925791873F01E2F69542805C3A3BC4B7FB0EF42512AF9;
defparam prom_inst_2.INIT_RAM_0B = 256'h3BA585A2F956AC3819B2F8492C06B7D6E2328EB646DD76D86E389910E9622675;
defparam prom_inst_2.INIT_RAM_0C = 256'h7BD5CDCE994B8DCC91447E3B3D93F090D80321CDA498335F7245597DFBDFECA9;
defparam prom_inst_2.INIT_RAM_0D = 256'h3389E264FC2C6D762EC80B9A0620ECA55E464A00023848DF6992737EC9A8895A;
defparam prom_inst_2.INIT_RAM_0E = 256'hB292E78677303749E7F58C888C91B72C8FE3034ABEB6B420047820240FAC3CCD;
defparam prom_inst_2.INIT_RAM_0F = 256'h11D3C4BD0A8D353F70512BD3F7EDA9D9B54BAE5B5C4C1FF57888105FE8E80940;
defparam prom_inst_2.INIT_RAM_10 = 256'h8B167EFFA3A95FCE2E66444837E9EAA792C39521912E5CCDAF71A1AACC9BEFC0;
defparam prom_inst_2.INIT_RAM_11 = 256'h3C1941AB79274100475564773A9840587D24464F858872370B31B99251CF71D5;
defparam prom_inst_2.INIT_RAM_12 = 256'h90F2E591E8724B577BD684008FAE5E05E47513FA1606FC9E7B83FCEB7D977341;
defparam prom_inst_2.INIT_RAM_13 = 256'h8B39ADE06C02CB8E8B9A0EAD37180BFD1D74FF7C9FA8F2F117B5C53DBCA8D6CE;
defparam prom_inst_2.INIT_RAM_14 = 256'hBC304FE0ADF236D1CEA8DFF7A4D33E53FB039FE272CC59EBDFDC26A76C067F92;
defparam prom_inst_2.INIT_RAM_15 = 256'h2AAFCB6C83DFB1DFEA865D8A67A0E0831DF99DB42EF7ECB9688BA6F3FFD183C6;
defparam prom_inst_2.INIT_RAM_16 = 256'h3D1D199FCF7A697FEF68716E6CA6E2746B379C6B444B9A9B576149BCD7D79A57;
defparam prom_inst_2.INIT_RAM_17 = 256'h60151AFFAD23F8A11DDC2E3EBA3D54A6D8E284CC3F7F476971E5907253D81052;
defparam prom_inst_2.INIT_RAM_18 = 256'hBC964F676E99F0749C4BAEF19DE71FE8F630FCC864048DB6188771CCBFE586FE;
defparam prom_inst_2.INIT_RAM_19 = 256'h310239E6EE5FD2CC954B02E449759885C2CEED90B7F73A83AB186AFA6609FE5E;
defparam prom_inst_2.INIT_RAM_1A = 256'hDF74411C8D64F5BC4097A54EFB1D6A83CEE0EBC7A9D37649EDAA427730D62293;
defparam prom_inst_2.INIT_RAM_1B = 256'hE5C8768AA9F76A444C083BDB48AB36CBA5B9E5938098A44E6E84779E9AB2AF54;
defparam prom_inst_2.INIT_RAM_1C = 256'h056E210CA388AD81A9C2265C928C2EC64FFE25367AF02B2974711F63C318EC47;
defparam prom_inst_2.INIT_RAM_1D = 256'hD2F76DBA26A3B2AF6B6ABCA2EAF37C241AE7A02D61FE5596A54B18A5828D52C4;
defparam prom_inst_2.INIT_RAM_1E = 256'h345F26E5BE0E371260F0E5BA71C3B1FE51B7C415CC31E9379BAC42DB049BACB9;
defparam prom_inst_2.INIT_RAM_1F = 256'h7913B36936A5B2BAE6296FDD4C5E191D52AB183049B52167679C085F36925F61;
defparam prom_inst_2.INIT_RAM_20 = 256'h298F827DE7320A1ED85764F919A8CCEABD0B7BECB90FC918F7F83B0B3B071A2E;
defparam prom_inst_2.INIT_RAM_21 = 256'h1602D76E351B7C4A694A185950D970005E0E26567E868BA471E26E06DF91AE8D;
defparam prom_inst_2.INIT_RAM_22 = 256'h5D9D4B6A02DFEA7A76356F31DBB0A920DAAE5FCF9ABFD04D3EDF1605F407E5F7;
defparam prom_inst_2.INIT_RAM_23 = 256'h5B67CB37CA4BE3297FE5D559AD37BA89826E732BA24CB9895555A90A3DB18D58;
defparam prom_inst_2.INIT_RAM_24 = 256'h2A3EAD8636FA1AFD71D418DA0F88B2BC573B6BE2EC5BFC7DD579602D0220ADF6;
defparam prom_inst_2.INIT_RAM_25 = 256'h5565E4E57506C8A6EDD27FCCD836BE09D492282D4F243DE08B153E175572D5FD;
defparam prom_inst_2.INIT_RAM_26 = 256'hDE0B6F19D5CB54E777F069E5DB5228D084E1267E3CBA86B28311D0C2CB47B1E7;
defparam prom_inst_2.INIT_RAM_27 = 256'h874CCA58CB2C75384997DDAAAAB72D47B6B141F4685A7A34AFA889F0C7D63EE8;
defparam prom_inst_2.INIT_RAM_28 = 256'h5C035ACF1B57D63F34FDD69AAB2D1658543D9ACB6E730A42C2CC6A4BF0FC7511;
defparam prom_inst_2.INIT_RAM_29 = 256'hA72DDE2F0605C88E3D5BCF176E602C8C14BA724F57E472A8E41542366803F68A;
defparam prom_inst_2.INIT_RAM_2A = 256'h134FA3EB419CBAD0194E189C63CBB67F79723010216548866427AD53821BFF37;
defparam prom_inst_2.INIT_RAM_2B = 256'h90E3AAB8FC6262B5B494060843B9DD78CCD78116995F2CC8048532E2B7BC3B6E;
defparam prom_inst_2.INIT_RAM_2C = 256'hE5D6572AE1389267F5BEDC1A1010419B3DA20171B2A28259AFD7A3DF5A0856EA;
defparam prom_inst_2.INIT_RAM_2D = 256'h08524A8293EA24A8BD8E551CE7D105315BA1A31601E74BE318CE37AB827299DF;
defparam prom_inst_2.INIT_RAM_2E = 256'hA3A032A84541CE042C8D3CCC84F5A2705C1DD30B964AF9CB1DA837C63F5BEFE5;
defparam prom_inst_2.INIT_RAM_2F = 256'hA11BC12F78CAE28DF6B77500D18DD95CFDC76CC0B41554E80B785F2BFC17E78D;
defparam prom_inst_2.INIT_RAM_30 = 256'h3DC2A7F1D611EB7C0DDEB070024B65E5EDB26D82BDF0038B36197F4F2E3F3DB5;
defparam prom_inst_2.INIT_RAM_31 = 256'hBE16B27F442066B1460936CD842FCE6BF9C3663E8E8C5E6990200717828E6124;
defparam prom_inst_2.INIT_RAM_32 = 256'h2F801C52FD1D4F8AFEECBB906548B6BCAC651AD16A77528D2634632CCD200E3F;
defparam prom_inst_2.INIT_RAM_33 = 256'h9C2C730AA08038FA7293F3C7F845B6125BBEA4B63EAEDB9C3A9EDF954CAC99EA;
defparam prom_inst_2.INIT_RAM_34 = 256'h3C460DB2A34D9866BF0071C2082BCA3B8C307E8115F62DF6E92199519D4ED6C8;
defparam prom_inst_2.INIT_RAM_35 = 256'h565C9CFBC4124596FBCACF328400E2AE5BD11B2A1420CE2F49116C244EE561EE;
defparam prom_inst_2.INIT_RAM_36 = 256'hAADA6215720FDF67B6F4879F629C37A90401C48FC639BAE5CEC63B29DD1EDAC6;
defparam prom_inst_2.INIT_RAM_37 = 256'h7878CA34EB24CC97ED122ECBA46DE716CC499B6AA6DB49A71D257A457036F6D3;
defparam prom_inst_2.INIT_RAM_38 = 256'hE5EB6D66458AABFCE4299A532CE2ACB28C08C95A396C4895596693454836E5DE;
defparam prom_inst_2.INIT_RAM_39 = 256'hF6DA4D1B88F5FB92B057150B2793297AC65E82DF2A0267F1ED242EDA258D2685;
defparam prom_inst_2.INIT_RAM_3A = 256'hC866049712349A072607FA892CBEE5F57C2634E38DE048B672A6B2E57DA12422;
defparam prom_inst_2.INIT_RAM_3B = 256'h11F45A6369DE6E74CB69343C3EB9C81DD227DA081C4C459D0009B1815B6CF760;
defparam prom_inst_2.INIT_RAM_3C = 256'h659B5F21378456D72D9922AB2CD26891EDC2993C3D3FE29DC098335123064D08;
defparam prom_inst_2.INIT_RAM_3D = 256'h5BC640A2F23F1F5635B5E959B8CEDB5491A4D3121EBF8C1F626B3B8A5D320B4D;
defparam prom_inst_2.INIT_RAM_3E = 256'h3057A71B278FB6DF98D0E504238E74E5E8C34FFFFC792639E08D3F48F56EA389;
defparam prom_inst_2.INIT_RAM_3F = 256'h2899BD57A5ADABC0EF19199B768961BDA7AEDEDC0E86900FF0E2CE38D86BFBD8;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[30:0],prom_inst_3_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 1;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'hCC36CE351B4DA9DAD799638B1E12042954965C3C1C9792E7BB6D3FFFE30D3E2E;
defparam prom_inst_3.INIT_RAM_01 = 256'h0CB4807FF1CB065F4C24402C1B7FD2B5BC06F6858190AC454A7A28D0909A403F;
defparam prom_inst_3.INIT_RAM_02 = 256'h5FC04B3D8B69FFFFCF24C7649A7E3AB5D422717D786B3CCBF70635A065F445EA;
defparam prom_inst_3.INIT_RAM_03 = 256'h79EEF9E06E5A8D8564D201FE18D9C7590B0DE9E5159CF136F15EF597B293C714;
defparam prom_inst_3.INIT_RAM_04 = 256'hC5826DF4BCA42A01C639D48D09A7FFFC71A7CF9E8391E9AE68C16AC9E0049059;
defparam prom_inst_3.INIT_RAM_05 = 256'h00000000000005F6D5D5FC28085AC72012C0E7F9749962A0BDE64F328072B713;
defparam prom_inst_3.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[30:0],prom_inst_4_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 1;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'hDC6F093738C0C3909FF80C7B9BAE67FB8807F8FFFFF8787B4DE386366497812F;
defparam prom_inst_4.INIT_RAM_01 = 256'h325C672528DF831E31838EF58FF07386455C8FF7000FF0FFFFF0F1F6996F1C64;
defparam prom_inst_4.INIT_RAM_02 = 256'h3FC3DFB6D0F9D976A947E6BC630E287FFFE1FC7503B31FE7001FE0E01FE1E3F9;
defparam prom_inst_4.INIT_RAM_03 = 256'h007FE0007F87FC69B6E3E34D2A01AD9C4639CCC5FFDFB1EE0F064006003FC0C0;
defparam prom_inst_4.INIT_RAM_04 = 256'h4133008E00FFE000FF0FF097BC8F3969B6E0FA1C0C47FC2DFFF818389809800E;
defparam prom_inst_4.INIT_RAM_05 = 256'h000FCE08126E019E0001E1FFFE1FC12D2C1C5A9AE7F14918181C25B300C0E3CA;
defparam prom_inst_4.INIT_RAM_06 = 256'h61C3425C003C702FA4DC031C0003E3FFFC3F805A483316338FF22A3830718AA4;
defparam prom_inst_4.INIT_RAM_07 = 256'hBF09BE4D5CE235981E7FC7473FE7E67F187BF407FFE700B3F5F631C06F036470;
defparam prom_inst_4.INIT_RAM_08 = 256'hD7D8C3177E18E04AB6E39A403CFFCB9E7FCFCCFC7071F01FFFCE0167EBEC6380;
defparam prom_inst_4.INIT_RAM_09 = 256'hFC00C59FAFB18735FF0CA20D4788A5A0F9E3F33CFF9F99F1F800E0FFFF1802CF;
defparam prom_inst_4.INIT_RAM_0A = 256'h3F9F8FFFE0038B3F5F4D47729FF33A9896EFBE03F3C1E5F9FF3F33C73C3C03FF;
defparam prom_inst_4.INIT_RAM_0B = 256'hFCFCCFE30F033FFF010F167EBE3BC7C91FB1D02167A6B51FE7E03373FE7E6798;
defparam prom_inst_4.INIT_RAM_0C = 256'h9FFD73CFF9F99F8E07C1F800063E2CFD7C738F621FF3805424260BFECFF86CE7;
defparam prom_inst_4.INIT_RAM_0D = 256'hF361A7E33CFE679FF3F33F3E03E3F0001CFC59FAF8E79EB43DDDE928E612C9F9;
defparam prom_inst_4.INIT_RAM_0E = 256'h396040D2AD63373FC12686A7C703B3FA0B5CC039FFC6449CB3FFFC999BD50A55;
defparam prom_inst_4.INIT_RAM_0F = 256'hCFE00183324E6A85B6E37F3FC68D0D4FCE0B76A0B64F0071FF8C833967F00E71;
defparam prom_inst_4.INIT_RAM_10 = 256'hFE3B1DA59FC0216622C3CBB63F42671FD97FBA8FFC070196981C00E1FF198E52;
defparam prom_inst_4.INIT_RAM_11 = 256'h15000381FC73374B3F803F6474FD442B1433238FE5AFF587F82248AB38DC41C1;
defparam prom_inst_4.INIT_RAM_12 = 256'hE0D4274CE22C07C0F8676C967F00EFCCE4A24ED3C833F187965FB587F073F359;
defparam prom_inst_4.INIT_RAM_13 = 256'h2C5E5607C0C50015429A0FC1F06F992CFFFE19D92C826A1FCE193807CB2F2B07;
defparam prom_inst_4.INIT_RAM_14 = 256'hA3B33C0CD82CAE0783C0E0FD9A141F83E0CF3259FFFCCBB26855E85BEB901C07;
defparam prom_inst_4.INIT_RAM_15 = 256'hCF3D30329E0700D645FEA1458C3B5E4A9A573137199E5C765F1C251CDBBDA735;
defparam prom_inst_4.INIT_RAM_16 = 256'h9C639971E004082FD81C06A88BFD6E8176E2BCBDAD57D77E737DB71C9E36C076;
defparam prom_inst_4.INIT_RAM_17 = 256'hE64D0C2D38C6408046D9AEFCE06032238FCD630468656E84B6B22C38FD92F9D7;
defparam prom_inst_4.INIT_RAM_18 = 256'h6A06AF861BB64623F1FBB4DBD575C8F3C1C1DCFFC64AC1C83D4A4D732A794C33;
defparam prom_inst_4.INIT_RAM_19 = 256'h55947D35B5DF581CECCB714BE336DC2CAAB1F85C8F87B6874DCAFF1ED0DED92D;
defparam prom_inst_4.INIT_RAM_1A = 256'h6BAC6C5233A8FD9457F11A3131A71DF3C7C1E782930CD9083F1FA6EC74D431A4;
defparam prom_inst_4.INIT_RAM_1B = 256'hF1F98AAE15AB4DCADB516295580240E0664DC6E38E0FCCA1FECEBB18FC7F1E53;
defparam prom_inst_4.INIT_RAM_1C = 256'h828F7C883B6A9F2A6C64E5D19BB3169E399F179CCB6E62649ECF28DC6175F57F;
defparam prom_inst_4.INIT_RAM_1D = 256'h7F0B5D656A6593507680DA54D937EEB8F318DD31835C2F1996DCC4C93F9AAFE2;
defparam prom_inst_4.INIT_RAM_1E = 256'h52F31324F81677244877CFC0F38634A9B7B964CF1ECD3A790E946E132D398992;
defparam prom_inst_4.INIT_RAM_1F = 256'h86328C4CE1E62649B22A5D700DF1F781C8664841D96B8B72B5A9F4F532D64E26;
defparam prom_inst_4.INIT_RAM_20 = 256'hD106D3E207E41C9992CC4C9326F374E0741F4203C22600C92AFB070D25D3E9AD;
defparam prom_inst_4.INIT_RAM_21 = 256'h6DCC63218CE5A77B81B21D33259899260FB6018EC24BBB0739B319B229E1BF7D;
defparam prom_inst_4.INIT_RAM_22 = 256'hDA896ACAC6834B3FB9574D0785523E664B31324C1EE9EAB2C2AB8A0E2DD0B564;
defparam prom_inst_4.INIT_RAM_23 = 256'hCC87CE0540961978E67C0B06ECBE38E2AF8F2E60D923DA15737F5EDA29EFA01E;
defparam prom_inst_4.INIT_RAM_24 = 256'hDF7A6D388E5EB03935CC321DF965A42EB520F9C5DF198CC1B247B46AEB4C168F;
defparam prom_inst_4.INIT_RAM_25 = 256'hC91EE56B8BD4A429140DA1F3E05864F1F44010B79CDFDBE5BE29D983648F6A95;
defparam prom_inst_4.INIT_RAM_26 = 256'hF8F5660D923DCED779878420312FFB1C8BF0C63F1479E00F817020207C673306;
defparam prom_inst_4.INIT_RAM_27 = 256'h1E24A348F107CC1B247BBDAE511CED1611CA95ADE861CA7F82EDCF67F9CC51F8;
defparam prom_inst_4.INIT_RAM_28 = 256'h7ACDC7E17AA89F71E25B983648F7535D96DB97F2BBDB8A8B46C38BBE5966A0F3;
defparam prom_inst_4.INIT_RAM_29 = 256'h970E5C624AF6619A1493DC63C7AB306C91EEAEB9A6C57C12A08E9984CF8719F6;
defparam prom_inst_4.INIT_RAM_2A = 256'hC1613762FF832C399C76DD7F097309B1657B0B4F80F2ECA7853F35E7C941377C;
defparam prom_inst_4.INIT_RAM_2B = 256'h92B2D19FEACC94D53F042BA330CE8D680F2C99124477EE9F01C5D94F826D205F;
defparam prom_inst_4.INIT_RAM_2C = 256'h3857650FE1FCDFC1EFD60E1CDE17A086E31FF8FB7F8386A6910B997E128BB29F;
defparam prom_inst_4.INIT_RAM_2D = 256'h7D1CC9F835AECA0FCCEBDF702F0937DC3C208099DC39DBABE0864A0D948536FC;
defparam prom_inst_4.INIT_RAM_2E = 256'hFB8CC1D38FD496F00E5D940FEA14AF7E5E2B1E8678780573738C44895CA065CB;
defparam prom_inst_4.INIT_RAM_2F = 256'h39D12BCB19BAEDB602506DE038BB280F9669CE0F7E109274F0BC56ECCF009CA5;
defparam prom_inst_4.INIT_RAM_30 = 256'hC17DC3307090AA5A72A3D76D0F98D3C27176500CE32F6301596DF161E18BFB98;
defparam prom_inst_4.INIT_RAM_31 = 256'hC8A23DDB0267F8AC7F8CB202884428E6212494756537D81BC324E780B3ED2683;
defparam prom_inst_4.INIT_RAM_32 = 256'h7973783AFC9FA57F43600F1401E0B88921129217BCB928EA4A6FBC007DB7F5D2;
defparam prom_inst_4.INIT_RAM_33 = 256'h56767F007AFD93AB4EB69662F5BFF3F938493D06E50D3A8453F251D088BF3E00;
defparam prom_inst_4.INIT_RAM_34 = 256'h5F2598E2DD268FF010687FDCD30B6F9CA6C02A797B29DDB54DFE19CF83B0CA31;
defparam prom_inst_4.INIT_RAM_35 = 256'hBD4F22D9F6697153AA0403F032B1594A6622FB44F40027C315E1C0F645AAE659;
defparam prom_inst_4.INIT_RAM_36 = 256'hD3EC07B9E06FB905EADAE2B64C0D81F0FFD16674162FF56C9EFFF487CC7FD1D3;
defparam prom_inst_4.INIT_RAM_37 = 256'hB40050DDC716DC31EF446089D1B5C5EC141B81F1F3585411821A00C2F000C35F;
defparam prom_inst_4.INIT_RAM_38 = 256'h88F03B11BFAB3664F4B4EA62E6B0C716EE7BB6EDD1E7FBF3EAEEEBFE5695F0B3;
defparam prom_inst_4.INIT_RAM_39 = 256'h0251CFC2672036DF7C832182B996664F49E7374FCCF7EDDFA3CFF8078262DECC;
defparam prom_inst_4.INIT_RAM_3A = 256'h4F3FE01E1237200263E0364AC2F4B8F2D8BE3E33AF7C2373D9EDDBBB279FF00F;
defparam prom_inst_4.INIT_RAM_3B = 256'h67E4EEAA9E00003C36592DF5237029244086BFF7D9CF4544490032B9F3D33756;
defparam prom_inst_4.INIT_RAM_3C = 256'h1E3E12FECFC9DD453C007FF80FF29B49D2783246B90545B2BB6E2B31F75A7B66;
defparam prom_inst_4.INIT_RAM_3D = 256'h4B477848A79C6B4B9F03BA0A7800FFF0EF55E169C9F8BE787496A3FAD1391259;
defparam prom_inst_4.INIT_RAM_3E = 256'h9DD7C202E86F73DB17FAC3573E07749CF001FFE100CAAD29BBF8DB073CC4482F;
defparam prom_inst_4.INIT_RAM_3F = 256'h7A0CC12807839F6B72E71C33755B276FFBB0952ADFFBFFC3A37F82E7DBF31C87;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[30:0],prom_inst_5_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 1;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'h0AB38EDFF3EC837144BA54CAA84268F58FC71A0FF7612A5DB0080000068F8997;
defparam prom_inst_5.INIT_RAM_01 = 256'h0020001FFF50C2AE911D9E19309B0F1FCC1BBACAB89B8BDFEEC254B140100000;
defparam prom_inst_5.INIT_RAM_02 = 256'hBB092D32FFFFC03FF6AC3B7C64D9CAD4DDA1E34F62D5ACAC66653D7FDD848029;
defparam prom_inst_5.INIT_RAM_03 = 256'h08C74DFF76125A5BFFFF807FD127B6601B19AD1F8B886B6792443AE63F50C3FF;
defparam prom_inst_5.INIT_RAM_04 = 256'h95D4459EC0335BFEEC24B5B400FFFFFFEB612E1D5A992ED210A1DEB2668167AA;
defparam prom_inst_5.INIT_RAM_05 = 256'hAEB9BB8277EDE671D4E7EBFDD8496A6801FFFFFE2E3874DA85906C63FED39669;
defparam prom_inst_5.INIT_RAM_06 = 256'hE211A61CA7D0C8C40923E236DFC077FBB78802199BFFFC006226CC760F30E0BF;
defparam prom_inst_5.INIT_RAM_07 = 256'h9CCCC0F99FA27E0FC0731790E9AD27E11E29FFF76F10047370FE7F3B389E48A4;
defparam prom_inst_5.INIT_RAM_08 = 256'h03F9F8F9BD60E25BC0171FED737376F3BD74928484D5FFEED63FE8BCC1FCFC78;
defparam prom_inst_5.INIT_RAM_09 = 256'h037FBECC87F3E3BCC1C00A6279175C68DD5C10C574ECD31E68F4FFDD857FD573;
defparam prom_inst_5.INIT_RAM_0A = 256'h70C3FF760EFFBC338FE78E6B9E87065B0D25B60F94F86320FA940D5882E07FBB;
defparam prom_inst_5.INIT_RAM_0B = 256'h3F613B9E54A5FEEC1DFF74CF1FCF18AE589B78AA2D512E3A47D63D86F7483D3C;
defparam prom_inst_5.INIT_RAM_0C = 256'hDAEFD3E089670897E47BFDD83BFEE99A3F9E716F05ADD73B8D946A199BD5A2BF;
defparam prom_inst_5.INIT_RAM_0D = 256'h6935918638DA4D61E8A1B468E0D38973CE7D21247F3CE3CAB3521AE2399C4A6C;
defparam prom_inst_5.INIT_RAM_0E = 256'h3662B9DEB4B374CC77A5A587325E410B622702E79CFAC24061FFFCFDCA035306;
defparam prom_inst_5.INIT_RAM_0F = 256'h9F9FEB576112895D6CDC043C3F35F60674C565D311C705CF39EFE481C7EFFEBE;
defparam prom_inst_5.INIT_RAM_10 = 256'hE7D6120E3E3FE36FAC90B5E3CFA0EE4CF2BBE05C1E8687C307860B9E73D4C903;
defparam prom_inst_5.INIT_RAM_11 = 256'h0C8E2E79CF5F2418707FC3DE64DED2055ED24A937E8DBE0904BDA9DEF78E173C;
defparam prom_inst_5.INIT_RAM_12 = 256'h88480ABAC79E5CF39EA648F1C0FF57D083D69279FB4620279C24BD69019B6BE4;
defparam prom_inst_5.INIT_RAM_13 = 256'h354AA4673DD7DDA28F1CB9E73C0091C703FE36DF5A57383BD4563120AA108C36;
defparam prom_inst_5.INIT_RAM_14 = 256'hEB61073F8B55F7E8BE883D58EAEE8F6EADD99B8C0FFFF693EEA7F6C773FC2A40;
defparam prom_inst_5.INIT_RAM_15 = 256'h590080C132C206DFE2967F47565740E935D81ADD5B31307AA1234CD9989057FB;
defparam prom_inst_5.INIT_RAM_16 = 256'h81E31FE39E3C717FC499885BE94939DE95F08470637121B7BA0320794386C1E7;
defparam prom_inst_5.INIT_RAM_17 = 256'hA2643C23DA7F19EC8FB837F80D26D0E06BA9DD40FA734146E683C36E5426181D;
defparam prom_inst_5.INIT_RAM_18 = 256'hA22E162A44CC3F7F1A0F8FC7CE8BC776CB57EB8BFFF8C53ECFD9CE9ED517025C;
defparam prom_inst_5.INIT_RAM_19 = 256'h98B1A82344FCA4541BD80F0FE3E733EC5818227397AA47DD1D78BA87A8C9CEE6;
defparam prom_inst_5.INIT_RAM_1A = 256'hB5C7A3C7CB6F7B8E91FBC9883FB00F981FD2304915B61BABA73A7F14F4B44F86;
defparam prom_inst_5.INIT_RAM_1B = 256'hCCF740D1C3F9777E65877AEAA7F9A4B7F70004DE58A620A6AFF7D66B6F800ED2;
defparam prom_inst_5.INIT_RAM_1C = 256'h7CF62302BC5493A088A182DCB74FE3B54FFB496FEE08C385D0FC3321B0FAA6E4;
defparam prom_inst_5.INIT_RAM_1D = 256'h7E065B9576C42B826A8D24395E838ECEA82B3CA8DFF292DED80C7E3CD7F560E2;
defparam prom_inst_5.INIT_RAM_1E = 256'h83C3F8F580FFA8A4A9CE82E3DDB860CE50D25CF679715298BFE765BD80C0039B;
defparam prom_inst_5.INIT_RAM_1F = 256'hFF8B96010F1B8C199F8CB40F3BE43700530BBFF401F7642AB49192317FC7CB12;
defparam prom_inst_5.INIT_RAM_20 = 256'h1B0EE157FED72C123F34C71EF03385A719C7627802653DD009FDE62A1EBC4B6B;
defparam prom_inst_5.INIT_RAM_21 = 256'h1089F634B86B9EA7FDAE5824FE54300002071FD621D77B9939E4583E25AC4061;
defparam prom_inst_5.INIT_RAM_22 = 256'h51AB932BB777C4492E4D87B38FEE94B899D5C7FC1E188F6C3A1C849BAB9068F7;
defparam prom_inst_5.INIT_RAM_23 = 256'hD64527BA6805FB298726F2EF1E51E378EFD9680ECC08C187FE66F69A3EA7E165;
defparam prom_inst_5.INIT_RAM_24 = 256'hFCD25019C2E10B072D7FF3D86D14BBC92D6B034E3FB6D1F982BF038FFEC01106;
defparam prom_inst_5.INIT_RAM_25 = 256'h0D43F3FFD9D452C7482884F44B3C888563F74CA837FC68CC7F6D8444D860E39F;
defparam prom_inst_5.INIT_RAM_26 = 256'hFD3D0213CB09F1FF9BEAE91F6CB87CD18A56F6950A0167B841C49CB8FE9E0E64;
defparam prom_inst_5.INIT_RAM_27 = 256'hF4863F1DFAD20BCD622C7000335701BDAADB2B6A1A2FB9162000D74D1578A431;
defparam prom_inst_5.INIT_RAM_28 = 256'h881F76B690C4D9CFF5A4AA621CA87000274E1115274AC8FC5557E37BE7FC8576;
defparam prom_inst_5.INIT_RAM_29 = 256'hC4AEE7883FCB389E01382CB9BBF66E55909070004DFA256C8D612E8D99B62640;
defparam prom_inst_5.INIT_RAM_2A = 256'hBB8E2A17E708C4D6CEB98A43D9672A4377EC4A40ED75483F80A206D8D7A70111;
defparam prom_inst_5.INIT_RAM_2B = 256'h1FA9B8451F8A13DD74094DAA817203B30F78EB86EFDF66ABE72D401F03DA4BDB;
defparam prom_inst_5.INIT_RAM_2C = 256'h000A7E3C132A50A6AF8A3E024C50A212865E2043778CCC8DDFBCE95B1DA85C1E;
defparam prom_inst_5.INIT_RAM_2D = 256'h7ED15B824CEB0FF81A472114C29F75DB14C87AC4D11723D4764B8E9BBF67ADCD;
defparam prom_inst_5.INIT_RAM_2E = 256'h474BC66EFD38A7F6052907F0D7FFB91BD3D0CDFEC1DABA6497E3AD4879249C37;
defparam prom_inst_5.INIT_RAM_2F = 256'hE749434EAC4744DDFAA72A7BEBA901E0D39D4DF5E4D475235334A81D674B140E;
defparam prom_inst_5.INIT_RAM_30 = 256'hAB34DBF40A944D0D20D315C98A36DD41F75B83C0C162E7260A9BE1A85029D2F8;
defparam prom_inst_5.INIT_RAM_31 = 256'h75EF357B98E90251874CA305B678DB808663650F3EF3878CD818B071E2B2BC8E;
defparam prom_inst_5.INIT_RAM_32 = 256'h8CF440E64615954C523777256F5412C9F3ED7611D486D9A23A4387100BD36660;
defparam prom_inst_5.INIT_RAM_33 = 256'h0A23CE21441A3A2C6A15D5D89989D8C6D4A9D55D9FB9CD33AE49126F97C38613;
defparam prom_inst_5.INIT_RAM_34 = 256'h4EDBE2820F738E4817E108F8FE54445ECCFE75B5D53560E0756F3338ADEDED86;
defparam prom_inst_5.INIT_RAM_35 = 256'h5D408F18C92CFD45BF710CCF02325C328E5666B96600C30D1F91F36045ED4631;
defparam prom_inst_5.INIT_RAM_36 = 256'hA71E2C7764853E3A90B132D3C6711DA365086E080F6751731D09D6B61C0CF7D7;
defparam prom_inst_5.INIT_RAM_37 = 256'h33DCDD4BF6754254754694A11BA45A29B8623CAF6EB3C5FC5AA4558A654060D8;
defparam prom_inst_5.INIT_RAM_38 = 256'h9E860E9427B02864F3220B6005050948F54FF9223398C49B0B505BB851C30B42;
defparam prom_inst_5.INIT_RAM_39 = 256'hBD8872265D20DA7C4C85A0D3C3E997DED61892974ABFF29C17318D3594FE9EA3;
defparam prom_inst_5.INIT_RAM_3A = 256'hA383B2ECFA6F95C14BC18D2E78EE3B6F230DA39DBE86250A747FF2FA1DE39B6B;
defparam prom_inst_5.INIT_RAM_3B = 256'h8BFFF5A7C767B4E7608FCEDB7A92B48EF68E25E4CC0C175E81B8CA26EDFFD73D;
defparam prom_inst_5.INIT_RAM_3C = 256'hB6EF28BF55FF79AD8CC7687DE3C74705A57DD3473426C3981E40354E51C59439;
defparam prom_inst_5.INIT_RAM_3D = 256'hFABAE88CE152501EAA010C5439CE5896A4D515155F3E6C8462AD10FE7777BC68;
defparam prom_inst_5.INIT_RAM_3E = 256'hC34FA542E65B9BD6C9C55F20BC027278538C9042D9A9082702389388DBCED58D;
defparam prom_inst_5.INIT_RAM_3F = 256'hF5B295BB3354707CD95CC7F45388B653F80000664E0734F63E033763CDBEA29E;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[30:0],prom_inst_6_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_6.READ_MODE = 1'b0;
defparam prom_inst_6.BIT_WIDTH = 1;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'h89933A65A54D4B40F75856E59A654F12A71B607D100002978C0E61278A60629C;
defparam prom_inst_6.INIT_RAM_01 = 256'hFC0DCE85E03204E576EA76907E26B813C6F56ACACE34F705E0000B641C0CE2A7;
defparam prom_inst_6.INIT_RAM_02 = 256'h7F8020777E198CFAF53EFE1563EA6649199C7E6C579404311C6AEE7C7FC00604;
defparam prom_inst_6.INIT_RAM_03 = 256'h70E8CA7EFF00428F7F13CDA05DF5A00A1F2BACE075914ADBE8849B6238550303;
defparam prom_inst_6.INIT_RAM_04 = 256'hFC680908E0D393F1FE00E7DC7F3350E030579B79FDAD484FFD01F128E71F3B6C;
defparam prom_inst_6.INIT_RAM_05 = 256'h52F607C76952978DC95C2643FC0001F87E64EC290AF2D5143E5295628CC3BFBE;
defparam prom_inst_6.INIT_RAM_06 = 256'h9BC53E98A0EC8787D00E22BEB2B7E99F0601F940E47DD5C71D80F1834ED92DF9;
defparam prom_inst_6.INIT_RAM_07 = 256'h319E1821359997E7DF7BF5D0DA1FF09C857046707E03CC81C8EB32B8FAA7F2A5;
defparam prom_inst_6.INIT_RAM_08 = 256'h071AFE3656186B49FC14CF84366A49FF9C0F3A508A64BB1FDF0CE0038184BE2F;
defparam prom_inst_6.INIT_RAM_09 = 256'h83AA9D8E1C761F3C7BAE4FA5D8529F01127D753DCCAF2E8D4AAACC7E0FD25587;
defparam prom_inst_6.INIT_RAM_0A = 256'hA937CD7EC06D231C30E1C48F9E3E53714D5A14A6E962307BA04D8CD394A53307;
defparam prom_inst_6.INIT_RAM_0B = 256'hAEE92A83519B33F9E0C45E38E3F91D5E57C03F8B2F4880A5256A5414702E8EC5;
defparam prom_inst_6.INIT_RAM_0C = 256'hA51125084338F585B1007A07C3E5BC73C7FD24C65BFBBEDBBCD45BC1B6FEC54A;
defparam prom_inst_6.INIT_RAM_0D = 256'h380F4BBD485160A453217B096710F46339BF56A7F96751A7F8A489AF0E780DEE;
defparam prom_inst_6.INIT_RAM_0E = 256'h7515F0449A0BD41A8E7007B8CA6A361A4463F386717A8D6FF2CF5AAF2A641F0E;
defparam prom_inst_6.INIT_RAM_0F = 256'h0B39F9C5FFCA168A7855EAB5157E996A28B9AC36D24FFFECFB918AC0058DFFC5;
defparam prom_inst_6.INIT_RAM_10 = 256'h956795FF96317965C71262E5256E5E6A79545A6ABA055824887E2B59FA48DAC0;
defparam prom_inst_6.INIT_RAM_11 = 256'hA1E16A67CC682BFF2CE8387CF6629445C67931D4E1E166BC480CB049FFF08FB3;
defparam prom_inst_6.INIT_RAM_12 = 256'h4792C0B4F783D8CE9E0453FE59E05F616903B4849F1C1DA85683ABEA022D60D3;
defparam prom_inst_6.INIT_RAM_13 = 256'h1EB3F3242E6D9408C82B019C3F98A400B192A481E596080BA2583F50E3355E4A;
defparam prom_inst_6.INIT_RAM_14 = 256'h0553B2DE8EB55718CE4300F17787A7B95AF787F9EBB081FAD12CB52894B19967;
defparam prom_inst_6.INIT_RAM_15 = 256'h05AFF271D4BF46049C9D0BBC2D1321E7B107169291BD5F3B1D620AEB7379114A;
defparam prom_inst_6.INIT_RAM_16 = 256'h0A192A6906D68D97C1195505972FB309A9C05FBC8F5300C6DC364D3866648821;
defparam prom_inst_6.INIT_RAM_17 = 256'hE8E6135A64B3B33F3B69D13D96533E54AF89632FD4CA787D6951AE0E1EB5256A;
defparam prom_inst_6.INIT_RAM_18 = 256'hADD74D87EACA0F299E6FE95EF0F81F9F8F3F118BCCA85763556081121C16BE01;
defparam prom_inst_6.INIT_RAM_19 = 256'h64E03CD4437F1911DE6D567ECFBF9D66AC3EA70A95F83AAEC95EA585B23C1F82;
defparam prom_inst_6.INIT_RAM_1A = 256'h05D4A715C7BDAB63FB6FFE6F84FF8B7A5B7D2E9E784D096EABB046946507331A;
defparam prom_inst_6.INIT_RAM_1B = 256'h839AC93E71214B77730A994F66E19685CB5A0CB56EBC112CC2D6DE9119DE8A9B;
defparam prom_inst_6.INIT_RAM_1C = 256'h2D2ABA958F25C01341A9E4472265620A71C76D1197B42691392A353A99BDB347;
defparam prom_inst_6.INIT_RAM_1D = 256'h781BC4DC6249000E9A613DE6BB3EEA2D0112B992D581A7F4571C458A4EFA9989;
defparam prom_inst_6.INIT_RAM_1E = 256'h2EB51238D9465242B815380532D6041938CCDDEAC4EB4C953BB9C7B1DCCD659E;
defparam prom_inst_6.INIT_RAM_1F = 256'h0EB12AE5D69396F48ABD5ABD048B667BC47B2AEB14E0C9A90FB543DB3B7877D7;
defparam prom_inst_6.INIT_RAM_20 = 256'h44A48D8AE932A6FFF030D3DF6495589BCDA254A78CA6B085827A5CB965536B5E;
defparam prom_inst_6.INIT_RAM_21 = 256'hB960DC1865485F30A4D066834038D28DA17C97369F5729AA18AE0F95D1CC2105;
defparam prom_inst_6.INIT_RAM_22 = 256'hC22AA819356CE30D8291AE42C3D367DBE99E3D93CD923AD1A71B1254717EC489;
defparam prom_inst_6.INIT_RAM_23 = 256'h9C6B56968494BFFA2AAFAF6B65742075D1989CFF713C749CBB247CA34E3C8198;
defparam prom_inst_6.INIT_RAM_24 = 256'h86AE04CB38EF8EB15C36FFC6C4D34CF7C2B694DBA08E56079318E719564854A4;
defparam prom_inst_6.INIT_RAM_25 = 256'hB363B1B9AC5EE534F18F4DEDD67301CD6564CF3B25502AF1B77675BD3331F7FD;
defparam prom_inst_6.INIT_RAM_26 = 256'h28EA86BD33C7DF134D4DA5C9E36892A9043FAF2C9198C7F4568358685AEE8B1F;
defparam prom_inst_6.INIT_RAM_27 = 256'h51EC012421549FF4278EBEB69A8C6797C7A0C720B0E9AD910EA474F7ACD5089F;
defparam prom_inst_6.INIT_RAM_28 = 256'h422DED0548E004814D453CCE671EEF4D35094F6F8F0BD64D338E2541E6EE4DE3;
defparam prom_inst_6.INIT_RAM_29 = 256'hADBDE7947A76356A9B63E3CFF8387272B47F96353DEEDB3018904AB7AEF13750;
defparam prom_inst_6.INIT_RAM_2A = 256'hE2CFA1897B648FF7E2E0B335356B58AA97B6927D60E3BB7A3BFABE60795B3F6C;
defparam prom_inst_6.INIT_RAM_2B = 256'h10493307CEF068E62701470E6F168DEA4E43AEE187CE3EDA8396CF9640455D81;
defparam prom_inst_6.INIT_RAM_2C = 256'h1C4B25A6DFAAE41F96AC4D8403D8E592BA166CD4EE24E323C798DCF506311786;
defparam prom_inst_6.INIT_RAM_2D = 256'hA2D94FA9709450E502DB99FC250899A131006D7381B927A967951891CE638ACA;
defparam prom_inst_6.INIT_RAM_2E = 256'h93AEA3736F72EA53E3969F46815633F08DAF0F0ED8BB639848E88F53F725EE64;
defparam prom_inst_6.INIT_RAM_2F = 256'h5017CF1C36127BD74B066CAFCFBB1AC9F6A84FC387560F5AEC00289ABACF46A6;
defparam prom_inst_6.INIT_RAM_30 = 256'h7FF359C56C50271D5F25EEC5EF16ADA6B7B348D26EA7F8781B1598C59F8FCE8F;
defparam prom_inst_6.INIT_RAM_31 = 256'hFD819D3B1E434C98FA04EE37C78003F5C0CA1378E0FE95CC5D4FF0F1CD577B34;
defparam prom_inst_6.INIT_RAM_32 = 256'h8AFFC3E67A8241A9EB2A1A223C1B0E445B9C3C175700607A98D968B477BFE1E3;
defparam prom_inst_6.INIT_RAM_33 = 256'h80C9AE26B57F87D43E18BD57599EC7B5CF6B1C127E7107CA64418203EFF6E886;
defparam prom_inst_6.INIT_RAM_34 = 256'h5A64AE99E996C5A3D4FF0FAE04B4C60F614661C388BD1C8BBAE5E55062D0669A;
defparam prom_inst_6.INIT_RAM_35 = 256'hC1C1325D6A78A4F58E6D447529FE1E7B81893B0D9B099CD407B31D88E02335E0;
defparam prom_inst_6.INIT_RAM_36 = 256'h5277AB40602CB8EB74C035BA78D2A96257FC3D69FDD2E62DF28141C1A98E38C9;
defparam prom_inst_6.INIT_RAM_37 = 256'hAF745C95488F5261C720B875520C118EC6D3F52CC1C389C60F8283BA46C156EF;
defparam prom_inst_6.INIT_RAM_38 = 256'h16F0942B180CCAAA307EA37FEDE05D5FEE5E92B35CCBA259971713816D833C6F;
defparam prom_inst_6.INIT_RAM_39 = 256'hF1DC4E0B477D9052642A2D3065FD4EAA9456F87723665CEB14B02A633C6E2705;
defparam prom_inst_6.INIT_RAM_3A = 256'hE526D29B8E389C3BB714522C82ADB98F59FAC0CE6B1B9E6CF8EE52C5D4FEB284;
defparam prom_inst_6.INIT_RAM_3B = 256'hEF0C00F7A5A05B67387138C71CC0F4C3AAA739F8D6F58908CEA67BA326133E3B;
defparam prom_inst_6.INIT_RAM_3C = 256'h90195904BA78D24C669B94CCE2E27076F4788D07EB00509897EB4BBE973A1D8B;
defparam prom_inst_6.INIT_RAM_3D = 256'h91B44D64C3552F071778D8D16DFBB39B8DC4E0ADAFFC1411B426F8F61FD7C39A;
defparam prom_inst_6.INIT_RAM_3E = 256'hBF05F3375369268B88CECCE1FF860F67EC8A100007863838A6B2692A5E158198;
defparam prom_inst_6.INIT_RAM_3F = 256'h5FDC162F3D370258A6D14A5141DACA323C90F2ABD7142FF00F0CF036723F7E79;

pROM prom_inst_7 (
    .DO({prom_inst_7_dout_w[30:0],prom_inst_7_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_7.READ_MODE = 1'b0;
defparam prom_inst_7.BIT_WIDTH = 1;
defparam prom_inst_7.RESET_MODE = "SYNC";
defparam prom_inst_7.INIT_RAM_00 = 256'h3007300615B9D373DCFF10B90D8B624EF089C5B814BAE95054285FE01C11C035;
defparam prom_inst_7.INIT_RAM_01 = 256'hDD217F80018C786A4677664C9727A4451B1FD391E92DB2A1D0B6F29010108000;
defparam prom_inst_7.INIT_RAM_02 = 256'hFA143D82DA42FF000F38F8515E635C11D81BCC5736B4546FB140F4D74E9268DE;
defparam prom_inst_7.INIT_RAM_03 = 256'h4577FB52FC1F3880568400001EE1F990DAC0FFCE558D9A6C6C83506D0CEC27DB;
defparam prom_inst_7.INIT_RAM_04 = 256'hB50CC7CF18A6389FC1FBE985AD0800007DC7F07F52A00AC9B88FB6B4DBB0B21A;
defparam prom_inst_7.INIT_RAM_05 = 256'h0000000000000C2F16969678E051B7C6A49DD0064231BB3B37F893884A4C94B9;
defparam prom_inst_7.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_8 (
    .DO({prom_inst_8_dout_w[30:0],prom_inst_8_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_8.READ_MODE = 1'b0;
defparam prom_inst_8.BIT_WIDTH = 1;
defparam prom_inst_8.RESET_MODE = "SYNC";
defparam prom_inst_8.INIT_RAM_00 = 256'h602F0237C7070121580007813031E0007FF807FFFFFF8783891C03E1B0B783D3;
defparam prom_inst_8.INIT_RAM_01 = 256'h242068A2505F923FCE0C0C37C0000C0220638000FFF00FFFFFFF0E07121017C3;
defparam prom_inst_8.INIT_RAM_02 = 256'hFFFC2038D801C070F0FFD03F9C1036AD0000006D30CF0000FFE01FFFFFFE1C1E;
defparam prom_inst_8.INIT_RAM_03 = 256'hFF801FFFFFF80071A603C1A1B1FFAD1FB801DBF9000041DD99BE0001FFC03FFF;
defparam prom_inst_8.INIT_RAM_04 = 256'h7BF00081FF001FFFFFF000E7DC0FBA21211F8F1FF007CFF00007E07855780001;
defparam prom_inst_8.INIT_RAM_05 = 256'h01FE0E31F7E00181FE001E01FFE001CFBC1F7C43400FB41FE01FCF16003FFCDD;
defparam prom_inst_8.INIT_RAM_06 = 256'h81FE034403FF804C6FC00303FC001C03FFC0039F783DFA82C00DEE3FC07FDC30;
defparam prom_inst_8.INIT_RAM_07 = 256'h7FFDF2764135B36001F83E8967E7E607E0000FF80000073AF424183A9FFCD47F;
defparam prom_inst_8.INIT_RAM_08 = 256'hD09060FBFFFD739C85DA1E0003F03C02CFCFCC0F80000FE000000E75E8483075;
defparam prom_inst_8.INIT_RAM_09 = 256'h0000F9D7A120C0F9FFCE16A92AED8E6007E018059F9F981E18001F0000001CEB;
defparam prom_inst_8.INIT_RAM_0A = 256'h7FFFF0000003F3AF424DC0FC9FCDBA507893B3400FC0318B3F3F30383C3C3C00;
defparam prom_inst_8.INIT_RAM_0B = 256'hFCFCC003FFFFC000010FE75E84BAC0CD1FCC5AB08DF606801FE053167E7E6060;
defparam prom_inst_8.INIT_RAM_0C = 256'h7FFC7E59F9F9800FFE3E0000063FCEBD0975810A1EF0B96327896B013FF8AE2C;
defparam prom_inst_8.INIT_RAM_0D = 256'hEB04901CFFFCFCB3F3F3003DFC1C00001CFF9D7A12EB82543DDEFC4602BC1406;
defparam prom_inst_8.INIT_RAM_0E = 256'h38E50B64A6B8F0F839C07667C70393FC073F0039FFF87EFC263FFB9E1A1CE48C;
defparam prom_inst_8.INIT_RAM_0F = 256'h98E0007C31C9293445A0F0F03700ECCFCE090B6F81C00071FFF0F5F84C7001FE;
defparam prom_inst_8.INIT_RAM_10 = 256'hFFC3D7A131C03F3821CE374AC8E1E0E03E64799FFC07FE0D87FC00E1FFE1EBD0;
defparam prom_inst_8.INIT_RAM_11 = 256'h66000381FF83A74263805D7873D70BF7D330E04039C873BFF83524583F3C01C1;
defparam prom_inst_8.INIT_RAM_12 = 256'hE0BDC132CB300700FF874C84C70045F0E3B222424D7070006790F3FFF00FACBC;
defparam prom_inst_8.INIT_RAM_13 = 256'h3043CFFFC08C8693AAD20E01FF8ED9098E00B3E1E3D454025EF8F8000C21E7FF;
defparam prom_inst_8.INIT_RAM_14 = 256'hF470FC00E0879DFF83C35566B3441C03FF0DB2131C01AFC3E667CDE1B671FC00;
defparam prom_inst_8.INIT_RAM_15 = 256'h6FC2000171F8061F81099F3C2F3C678B23F7C6F7E61F9C5C00F88D37C77F7253;
defparam prom_inst_8.INIT_RAM_16 = 256'h83FCEC400FFA6810C7F0023F02131E75097CCF3EC8BCF80F8C7E3FA801F93A56;
defparam prom_inst_8.INIT_RAM_17 = 256'h07B1C16D07D8630021D9D1FE1FE0363C142300F242198CF92680291F01FCE696;
defparam prom_inst_8.INIT_RAM_18 = 256'h45D61EF81C47C4FB8F824B037331764DBFC1F4C03006002A54F38985F7FA023C;
defparam prom_inst_8.INIT_RAM_19 = 256'hC6E7A9D9CBC061E0F00C05FF1FA23B56E65E90D87F87EF00E1467FFF6DE71236;
defparam prom_inst_8.INIT_RAM_1A = 256'h0F9C7115DFCF5626BE017BC1C038E89E3FB451878FE1D2E0FF1F9BE346CCC16D;
defparam prom_inst_8.INIT_RAM_1B = 256'hF1FFDD9CDF9B8F6C679E2CD9D99ADB038473E93C7F4F42FC01D406D9FC7EEBCE;
defparam prom_inst_8.INIT_RAM_1C = 256'hD1D228B83DCC4625BAFD00B7E2E7CF1FC6DEA81F0D99B7DD9F40CF9783A6C03F;
defparam prom_inst_8.INIT_RAM_1D = 256'h7D31ADC3B9BD1AE07BDC884B74CDA7AAAFA94E3E0D92F01E1B336FBB3E8EA5F9;
defparam prom_inst_8.INIT_RAM_1E = 256'h65CDBEECFC7E0E439B958040F5BDF096EC3A4F9AFFA2FC61F30F301C36E6DF76;
defparam prom_inst_8.INIT_RAM_1F = 256'h87BEF070CF9B7DD9B8AD63CFFBEB7E81C007402D498D6A9719D438C6031CF038;
defparam prom_inst_8.INIT_RAM_20 = 256'h9711E3CB0760E0E1DE36FBB33177EAFFF27CF283805290129CB58A60C22871C9;
defparam prom_inst_8.INIT_RAM_21 = 256'h09F84A8AFFCDC65381F3E1C3BC6DF76623E84CD106446507B5B2200512F0A543;
defparam prom_inst_8.INIT_RAM_22 = 256'h7454841616A81B0190938E57814FC38778DBEECC4525216086E8840F7BA2420A;
defparam prom_inst_8.INIT_RAM_23 = 256'h69075606FEA6C4CD47D3F92B4BA03F3B180FDF80E63C111E59F379D8A5BABC1E;
defparam prom_inst_8.INIT_RAM_24 = 256'h6CCB3F9D0F9ED030B91D89912BD933C3DDF0F7A63015AF01CC78227CBB4D7FF6;
defparam prom_inst_8.INIT_RAM_25 = 256'h31E0ADB2DEA98E260CAF61FF675B13DF523FE070AD3FF4F660309E0398F046F9;
defparam prom_inst_8.INIT_RAM_26 = 256'h80E0780E63C15F65DA56A0C4277783DFC7B621A07D07CE85628FED77C064BC07;
defparam prom_inst_8.INIT_RAM_27 = 256'h8CE32EAF01D1F01CC7829ECB3A2662D85CA3E64AB0EC4092D98992DC61C3CCAF;
defparam prom_inst_8.INIT_RAM_28 = 256'h6C3C1488E4666BDE02CFE0398F053D967AE93CA1A2DDECD024D88AA2EC783F49;
defparam prom_inst_8.INIT_RAM_29 = 256'h136274C80CC5A72FB44C193C0697C0731E0A732E69C0F88C6080D16647B11D74;
defparam prom_inst_8.INIT_RAM_2A = 256'hC3643EE8E830FAB1E7876355655A23B679C18C702BB9F63806CCFD6C24C9A577;
defparam prom_inst_8.INIT_RAM_2B = 256'h1CC2594FE497DE3A0064FEA3CF00F0A8027D2DFC7BA600E05773EC70034888BF;
defparam prom_inst_8.INIT_RAM_2C = 256'h658FB1F021E7BE9FFDAE54E920DCFA071C1FE2C8B4A7E0D8FF5F4180BEE7D8E0;
defparam prom_inst_8.INIT_RAM_2D = 256'hFA588E02CE1F63F07C1015CFE281EDEA01B0C1DE2007EC5A9B4DFDB1FB4F8701;
defparam prom_inst_8.INIT_RAM_2E = 256'hE79C21E354FD1805983EC7F0999D2B01C56013AA835B6E7C0383B97B6F4C9B73;
defparam prom_inst_8.INIT_RAM_2F = 256'h3E1F5FE4D5E71BC738D6700B107D8FF1713B1F00ED9F777A06F286F00F009766;
defparam prom_inst_8.INIT_RAM_30 = 256'h19E8CFC07F22A79F3B0A8F8D65ACE01420FB1FF3E1D89D009280EAF20DAF1BE0;
defparam prom_inst_8.INIT_RAM_31 = 256'hC2735FCC13F7F81214015C814B96E1B47CB6F3A2E322101FC1409F81B2FDDEDC;
defparam prom_inst_8.INIT_RAM_32 = 256'hF4172C27BC999707800FFB4AF54FE702C4D4FD28E3EDE7454644200FFA0A7C4C;
defparam prom_inst_8.INIT_RAM_33 = 256'h3098003FE851B28CCEF5E5EF20E01DE3B9CA80DB55129CF2F85BCE8E98C8001F;
defparam prom_inst_8.INIT_RAM_34 = 256'hE7CBFD3A41F8700FF15CD6B2DC46E6D50C402CF528505B274C2F78649427FC9D;
defparam prom_inst_8.INIT_RAM_35 = 256'h06B9CC19E1B7FAF093B9FC0FF30D74241DC1EC3A69FFB93E473F992B0D0B34CF;
defparam prom_inst_8.INIT_RAM_36 = 256'hE04634B4C2412FAF5567F5E03773FE0FFFA9098A33CF68818600B5836602BCD0;
defparam prom_inst_8.INIT_RAM_37 = 256'h1801F63F33773A98513D51C0A2CFEBC0E6E7FC0FF0AE8761C3E312C316015115;
defparam prom_inst_8.INIT_RAM_38 = 256'hF60838DF8DD25F43E19CD40BF34070435780239BE060000FE40E27D4959A45A8;
defparam prom_inst_8.INIT_RAM_39 = 256'h086F139D86C03A63A9D7E1F6322F6973266DADA7AF004733C0C007FF8618F0C3;
defparam prom_inst_8.INIT_RAM_3A = 256'h43001FFE155D16E2504031B37AE5C7E5DFCC465BE3AA69ED1E028E67A1800FFF;
defparam prom_inst_8.INIT_RAM_3B = 256'hF819399C86007FFC278961F7818031557F9140048B7934A77F850C027C0D9CCF;
defparam prom_inst_8.INIT_RAM_3C = 256'h2D5A1433F03273390C00FFF80260186ED10066434CD5767355AEE994A67E63A0;
defparam prom_inst_8.INIT_RAM_3D = 256'hC7011DC71C720665E0F4E6721801FFF061B856639A00C5F9F5F0CB05DF516A79;
defparam prom_inst_8.INIT_RAM_3E = 256'hF6D83DB5C448602731FCB1CBC1E9CC6C3003FFE0F05F8EF64E0098F5B67C7192;
defparam prom_inst_8.INIT_RAM_3F = 256'h98C0FF6142445AC95CC9C520C58D3C280023F4CF8FFFFFC0169B867828001FD7;

pROM prom_inst_9 (
    .DO({prom_inst_9_dout_w[30:0],prom_inst_9_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_9.READ_MODE = 1'b0;
defparam prom_inst_9.BIT_WIDTH = 1;
defparam prom_inst_9.RESET_MODE = "SYNC";
defparam prom_inst_9.INIT_RAM_00 = 256'hFF30ED1CF010FF0D226355D97F5115F991AAE4700047E99F1007FFFFF9DB4811;
defparam prom_inst_9.INIT_RAM_01 = 256'h801FFFFFF857A905F6C1FFF8EEB4AE0F951CE6A925A34500008FD334000FFFFF;
defparam prom_inst_9.INIT_RAM_02 = 256'h023F1E1500003FFFF2D8266CDDA1F30F15D889F0AE9F728D21A93B40011F8F2A;
defparam prom_inst_9.INIT_RAM_03 = 256'h8EB18400047E3C0E00007FFFEB5B56094EE1C9F2601AAA25D13C51CC8F398780;
defparam prom_inst_9.INIT_RAM_04 = 256'h74E5F76200564E0008FC781FFE0000FF18230C8C48E1C856388AFDC2D2EBB76B;
defparam prom_inst_9.INIT_RAM_05 = 256'hCD097BE6930B7687A8FDC80011F8F13FFC0001FF952722B197E070D0C1CC24F3;
defparam prom_inst_9.INIT_RAM_06 = 256'h5D98EE0599431BE2E6CA912DD2C0200024E7F888780000038F9A1A421BC3007D;
defparam prom_inst_9.INIT_RAM_07 = 256'h7E60F40748B52E000026C6DDAC2BD283AF32A00049CFF150F001FF0211387795;
defparam prom_inst_9.INIT_RAM_08 = 256'h0007F813AC60FAFB05B7BFEF5AC1D56AAEF0093CED7880009B8002A3C003FC0F;
defparam prom_inst_9.INIT_RAM_09 = 256'h368016BC000FE061A0C0038437A21F971D377A46F35072D10BFAC0011F00014F;
defparam prom_inst_9.INIT_RAM_0A = 256'h550900046D00ADF0801F81DF2C80C47C78FB3872551D5D0C826F05F380458002;
defparam prom_inst_9.INIT_RAM_0B = 256'hE5B12DCAFC680008DA015FC1003F07FDEA87EA618B4737298E7EE3B3DC52997E;
defparam prom_inst_9.INIT_RAM_0C = 256'hF06D8DF189CDD0E8A25C0011B402BF86007E0F4E5F9DDF11434E4CCB29EABCB1;
defparam prom_inst_9.INIT_RAM_0D = 256'hC53120789D4B66B133C884660284085B4783D71C00FC1ED0633032148B0C9167;
defparam prom_inst_9.INIT_RAM_0E = 256'hAD8CCF5F75FC765A83FA87008D6AD0F7200800B68F072E301FF80018AEF466F9;
defparam prom_inst_9.INIT_RAM_0F = 256'h7F801643761CF3591EFC08AE1694A6412843B85A2A18016D1E043C603FE00E4B;
defparam prom_inst_9.INIT_RAM_10 = 256'h7846F181FE0004CF4D9CC7439600CEC2A912DB3549D474242C7802DA3C0878C0;
defparam prom_inst_9.INIT_RAM_11 = 256'h2BF00B68F0DEE307F00009430598D54CCE9B97B14B510DA3E381DF4C80F005B4;
defparam prom_inst_9.INIT_RAM_12 = 256'h211F74A71BE016D1E1BDC60FC00082D26D1850B8F16BE088B2EECDBE5ABE93C4;
defparam prom_inst_9.INIT_RAM_13 = 256'h7B386657CE6B57161BE02DA3C37B8C3F0000948CC3987A914C67F0607F46A865;
defparam prom_inst_9.INIT_RAM_14 = 256'h4C7FB46209D06AF168FA3234DB192BC1CCF7807C00013B518F3955767FFE7067;
defparam prom_inst_9.INIT_RAM_15 = 256'h4D7B55BCACFCDD8FEA0867296756EAA46637538399EF0FF99F1B8F6EC2AD9835;
defparam prom_inst_9.INIT_RAM_16 = 256'h7E1C07C1D6F6A9B498E8E41C3E299A40F9B0833064EEB30F3BDF1FF73078F1B3;
defparam prom_inst_9.INIT_RAM_17 = 256'hED1C43E023BFF8782DACB732B1CE4BC5E0E8FDCF7E27438349BD661F779E27FC;
defparam prom_inst_9.INIT_RAM_18 = 256'h3EF491ECDA3C80FF63FF96009A29572BF390CFF87030CB1AB4D93DE71B7A48BE;
defparam prom_inst_9.INIT_RAM_19 = 256'hAAC1B8407DE92BD9A63900F0FCE0AE3D715D09D4E72776AA1C55D13751069142;
defparam prom_inst_9.INIT_RAM_1A = 256'h850DB2C5F0CDA380F3D257934472001FFE300AC7E2BA12CDC66CCDBC5AAE5A10;
defparam prom_inst_9.INIT_RAM_1B = 256'h72D323845FA7BEA1CC522F9CE7AA742718FC00E1C79C7A73456F974F8D42B1F7;
defparam prom_inst_9.INIT_RAM_1C = 256'h2B6DF2DCC561EAA868BE5528CFEB92C9CF54E84E31F8FF84B70610101434714F;
defparam prom_inst_9.INIT_RAM_1D = 256'h0015DF014BBF96E38946A3AD599EC3C0D87E2113DEADD09C67EF8E0248034440;
defparam prom_inst_9.INIT_RAM_1E = 256'h7FBFC7CC40F66286E91664BC2B294AF33D0337F7C97106EFBD5BA138FFC00079;
defparam prom_inst_9.INIT_RAM_1F = 256'hF57A84E2FF07FC781FEE66439B420380611AFE342572CB36F90BB9DF7ABF4271;
defparam prom_inst_9.INIT_RAM_20 = 256'hED83E66FEBF509D5FE0CC0FEFF5C33A7414AC2F8B1C7072D56FB3C37772A58B7;
defparam prom_inst_9.INIT_RAM_21 = 256'h0063E19CCF44A0DFD7EA13ABFC320FFFFDC4E35EBAA0EC79EE4B30301883C691;
defparam prom_inst_9.INIT_RAM_22 = 256'h0FBB576EB1018A4A6C2C8FCFD4BE238F844C3C03E1180EFDD1F5C878B1E4D2DF;
defparam prom_inst_9.INIT_RAM_23 = 256'h5D613694F9A1FC211D9C7057EAEC745749784711CD47007801E0FFC387CDB7D7;
defparam prom_inst_9.INIT_RAM_24 = 256'h03C00D08D95F9F3D9A71491313196174577ECA40B2F08FD86180007001C99F87;
defparam prom_inst_9.INIT_RAM_25 = 256'h733FF00007D0CAE9B95B0D8B2D99A2C10CFA63D4AC37058165E13BFC07E0E060;
defparam prom_inst_9.INIT_RAM_26 = 256'h9706E2F07507F00007D751E9ED9E075A6E3624B802534F58159DFB02CB83709C;
defparam prom_inst_9.INIT_RAM_27 = 256'h43CA97172E25CFC3BAE3F0000F80B21D09A9EA3B2BD783D27DB4FCE0726551FA;
defparam prom_inst_9.INIT_RAM_28 = 256'h0FBB5AD1265040165C4B361D1A67F0001F2F6493C1CF9CF295B62EAF8C104E98;
defparam prom_inst_9.INIT_RAM_29 = 256'h9559FE99509066B46228C658FFA0E930EC4FF0003DC4CDC8C1881D95B0012BC3;
defparam prom_inst_9.INIT_RAM_2A = 256'hBB5A237FB1B80B52F872922F7BAE6BE1FF41D6CE399CC00783557A40DE2D25AC;
defparam prom_inst_9.INIT_RAM_2B = 256'h11FCF6D10D64FCD2F20F7899B619541F92C5E743FE84DD921B6CC00F02683749;
defparam prom_inst_9.INIT_RAM_2C = 256'h1BF9FE3C3ED9F44A5D0B806A11F239965C3F2331D358B387FD085B3D5559DC1E;
defparam prom_inst_9.INIT_RAM_2D = 256'hF43FC8FE5018FFF85DF09B1D0957F08B4072BFEBD95843312B8C288FFA171BCE;
defparam prom_inst_9.INIT_RAM_2E = 256'h29FA083FE8626F0DCA18FFF06D54939B0A96229055A189AF1C64B4FF78AD501F;
defparam prom_inst_9.INIT_RAM_2F = 256'h48E06448E1DA9C7FD043678ED398FFE0BB16EAB4313C2F134EC2E618992EA870;
defparam prom_inst_9.INIT_RAM_30 = 256'h329DCA77C6ADA1390D0F97A7D5B1C5A8BB387FC1645DD1A2D26B543A3B84C6F6;
defparam prom_inst_9.INIT_RAM_31 = 256'h7390C1A82DBB523A1FBA0AC508871F4F2960E1DF8E007F8068F6C59BD9C562E6;
defparam prom_inst_9.INIT_RAM_32 = 256'hB084DA090280164379564043F5DF2B809F28DE8E82DE3D9F67307F0A34212B24;
defparam prom_inst_9.INIT_RAM_33 = 256'h16603E2EEC719675A194F946EB0A2973280BA7611C37FC0D03C72400D6407E02;
defparam prom_inst_9.INIT_RAM_34 = 256'h49C77B01D7F07E56EA90150B667DA6C31A99870BF3F66F535A565902A6E3F600;
defparam prom_inst_9.INIT_RAM_35 = 256'hF7336712D31CF98390F0FC90AED805F4D6AD3A7D53F0E52E3625AF6E2E70B205;
defparam prom_inst_9.INIT_RAM_36 = 256'h258F66675FDAEE2FA4708496A7F0FC642D248E63B8196505B7D79ED777E30EDA;
defparam prom_inst_9.INIT_RAM_37 = 256'h5A42E1CBCB7B9E79AD9800C177612CA457E1FDBC90531B2B70129F9329C1FDCB;
defparam prom_inst_9.INIT_RAM_38 = 256'h8438E0E6B48F55C95159AA90040531832CCFFCA04167C47C7A5F3E063A474C7B;
defparam prom_inst_9.INIT_RAM_39 = 256'hFD69A1389D3DC3996A75130A3A93BAC2AA226301799FF90932CF8CF187E45715;
defparam prom_inst_9.INIT_RAM_3A = 256'hE83FB1DC37AAAFD927A20E34B5E1CED1015AE22F86644622723FE704341F98F3;
defparam prom_inst_9.INIT_RAM_3B = 256'h98FFF9C7D01FF3F722D47B625754B8EB6A67301590673FB92A2D0C58E47FDBEC;
defparam prom_inst_9.INIT_RAM_3C = 256'h537431AF33FFFDC4A03FE71CB71235795D97E394DF408B738DF1DE3ABEA518D3;
defparam prom_inst_9.INIT_RAM_3D = 256'hBB316CB2A29862CE6600882D603FC68B9E63D4A6B6238F29B612EA58FE9726B0;
defparam prom_inst_9.INIT_RAM_3E = 256'h94D1E64EBC5803518159981AD4011816C07F8C30E8C6AFA485DF1CD36A040BAC;
defparam prom_inst_9.INIT_RAM_3F = 256'h737CE6C5A928BC990BAB4DE2F2B131A7200004AEF9FF0E5D8C7692DE649F3B24;

pROM prom_inst_10 (
    .DO({prom_inst_10_dout_w[30:0],prom_inst_10_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_10.READ_MODE = 1'b0;
defparam prom_inst_10.BIT_WIDTH = 1;
defparam prom_inst_10.RESET_MODE = "SYNC";
defparam prom_inst_10.INIT_RAM_00 = 256'hCD5F82BDFCD18D952A0747968C84ABA0256274B640000956F3FE14F41920FCBD;
defparam prom_inst_10.INIT_RAM_01 = 256'h03FC382CDF356976B1CC7B0BB740BAD2A59265DF8AC6D96940001695E3FC19E3;
defparam prom_inst_10.INIT_RAM_02 = 256'h80007F4A01F861830C2E2D55E073F43FCB2898E6D6D24231158CB2A6800031CF;
defparam prom_inst_10.INIT_RAM_03 = 256'h573034E500008F4500F014D6BE08F32EFFCCC8131BC1E3024449F6572B99A54E;
defparam prom_inst_10.INIT_RAM_04 = 256'hAE06C46CAF600ECA00011FCA00F1098F8FA542E000319059BB28A6095404DC26;
defparam prom_inst_10.INIT_RAM_05 = 256'hC4F818CA876D94C01661A87C0003F1D401E2099BC65D15E43C6325D301F9A388;
defparam prom_inst_10.INIT_RAM_06 = 256'hD5A9B2DF8136ACF3447E4854DCCB01E8F805C2981BFE9B7F46DEB859133E4B6A;
defparam prom_inst_10.INIT_RAM_07 = 256'h182ACF01BAA2F25F88E182D36F01268D9999E79FF00BB73037EDB1F867EFF163;
defparam prom_inst_10.INIT_RAM_08 = 256'hFF2337CAAE073A0D30193B113E5279D57513BA5EF3B03C3FC014F6607F993DC2;
defparam prom_inst_10.INIT_RAM_09 = 256'hFC45F681FC07FADEC880FCB6146489FB5A623EAF1289BA31F341703E30200940;
defparam prom_inst_10.INIT_RAM_0A = 256'hCFF00F01FF9C2D03F001A0A2F8E37BA0F593C662DA08AC0E7AFE71E3E722C37F;
defparam prom_inst_10.INIT_RAM_0B = 256'hCBD1B4139E703FF9FF234207E001FA0BD011D7399C6E5A04CE11A72A8E9BABC1;
defparam prom_inst_10.INIT_RAM_0C = 256'hBD4564CD9843D2DE4E2785FFFE4E840FC003CA653533ACB7E898EE0BF5981FBF;
defparam prom_inst_10.INIT_RAM_0D = 256'h362F69C771E75617626155BC98BF03E0FD929E6002C4AC8091A638980F0904F3;
defparam prom_inst_10.INIT_RAM_0E = 256'hF873E578F4E8F38EE3C16C375B8F6B7132BC0C01FB293CE00588D841F0D6AFF0;
defparam prom_inst_10.INIT_RAM_0F = 256'h16057671938BA2F3ACA0E4DDFFF71F0E36FE16E032700003EE2EF9C00B0168CB;
defparam prom_inst_10.INIT_RAM_10 = 256'hAA6C73FFAC472FA1A00B74F6107C433B802019EB4248ADC0608058C7D54D39C0;
defparam prom_inst_10.INIT_RAM_11 = 256'h4000731F9698E7FF589A4B7A0C8CE769FB1105775B15F0446E2B5B80A600000F;
defparam prom_inst_10.INIT_RAM_12 = 256'hB8456E903C01C63F2CF5CFFEB109B56E1E1BD8D6A66A16EE7B39F33603DCB741;
defparam prom_inst_10.INIT_RAM_13 = 256'h24E7485FA29D0D99D2E6087E59FB9FFD601372DF78D0ACADBF9C29DC6DC53E9D;
defparam prom_inst_10.INIT_RAM_14 = 256'h82E9A78B1D9A8885E8F90BDA684D8EA0C34780061E6EE5A15A7666895B7CD3C8;
defparam prom_inst_10.INIT_RAM_15 = 256'h9D15638631CB4E98C1E8F733D73257A62B119F3180333034F7DFC4902BBCA9A8;
defparam prom_inst_10.INIT_RAM_16 = 256'hA3AE0BCC23DB0E2A5390CF4A8369D989F68433732BAB1D81CA72CE3D8D9F1C0F;
defparam prom_inst_10.INIT_RAM_17 = 256'h2C781C19A7DD8D9C918E6A2E57608C72A46B51B2AE97A687C9FB3841D23339B2;
defparam prom_inst_10.INIT_RAM_18 = 256'h2150840773ECFF56FBB3E57762001FD9EDC015308FCD9B59BAD34CF354194900;
defparam prom_inst_10.INIT_RAM_19 = 256'h00CD08890E7A681E787130B5644770C28DFF3611520029077FD15BB4EDDE8496;
defparam prom_inst_10.INIT_RAM_1A = 256'h1272D719F8FE5ECAB16A6C7173FF5A68488D847B283DADA02440611791306245;
defparam prom_inst_10.INIT_RAM_1B = 256'h3BCA610384FF15914AADF4A3885D4C4D59595C726B99E64E2B30999FD5F041FC;
defparam prom_inst_10.INIT_RAM_1C = 256'hB6F33A827784CAD70E877E9036EBE79F91764893CD4D6187B01A19BE527134C8;
defparam prom_inst_10.INIT_RAM_1D = 256'hC2ED491575F2329D6B16749D7B72DEC2FD1FB662D2B824840A853C644714A2F4;
defparam prom_inst_10.INIT_RAM_1E = 256'h69730E576ACAE468AFE60EB6D22CD5530E35478DBB3B652071BF297147C4E396;
defparam prom_inst_10.INIT_RAM_1F = 256'h87C6A9B1A78F8E6BF0E59329ABEC071685224FD44600FECBF134503823C9D2C1;
defparam prom_inst_10.INIT_RAM_20 = 256'hAE821546779F8195620FCE57C8106ED353CDFECD0A1552406FD5A144DA403EEF;
defparam prom_inst_10.INIT_RAM_21 = 256'h13D3F349B905F5ABD16F802A6407CE5A4CC8DBA7A3999953177714FE9ACBEDA6;
defparam prom_inst_10.INIT_RAM_22 = 256'hBF243DCB2B3B114C6A0AF7A790727DF5307E0225AEDB5C9E381D6426495B7916;
defparam prom_inst_10.INIT_RAM_23 = 256'hE060D53F5175F9D7C0B43B6C1401ABFF470AA6A0C0FC0A0E2DB6B13C70386E9C;
defparam prom_inst_10.INIT_RAM_24 = 256'h34F4C933C0C5156E17EF13746E8B5835A055137E2AE2D2CD90F806D41B6D66D8;
defparam prom_inst_10.INIT_RAM_25 = 256'h70E0061D49EB764701D31ED28BA0E4D8C41B2DDFC0BBC47A7A5368D170F010F2;
defparam prom_inst_10.INIT_RAM_26 = 256'hA9F02C85F0C0B3F49696C90E0370F7866ABB4F72BC4FE85B8967C772BEF909DF;
defparam prom_inst_10.INIT_RAM_27 = 256'h2C798DD6C05957FBE18061452D29B61806A4C12F1F813B6110D5D053121CE4F8;
defparam prom_inst_10.INIT_RAM_28 = 256'h5CC62381034D83D68D949631E302C7BE5A526C700D09C65D58EE9B9F4E114B82;
defparam prom_inst_10.INIT_RAM_29 = 256'h0DF86DDE1167FC020E18CEECADF4E5E98BF89F61A1489BC00049E7AF9779C7B8;
defparam prom_inst_10.INIT_RAM_2A = 256'h15F8B53F5D032C2B4480D1A41EBA85CA340792531FE6420342B33F8000B9DB5F;
defparam prom_inst_10.INIT_RAM_2B = 256'h1A8DFC000B00C6E9CBC241AC7330E4883EFA45E119250B867F976F8485667E00;
defparam prom_inst_10.INIT_RAM_2C = 256'hFC16E834EA3378004D718BF4CF90D200BFF1B2100049E90A2BDAE44CFE2C23CB;
defparam prom_inst_10.INIT_RAM_2D = 256'h6DF6B067F0FA6DC9D4ECE1033438038B8FD11DA8FE3B94201C3E8A762A55AFB9;
defparam prom_inst_10.INIT_RAM_2E = 256'h0DBED71779AF9BCFE1282D972999C20F2129EAF47631B505A603D241300F1A91;
defparam prom_inst_10.INIT_RAM_2F = 256'hD521053DB16C97846C5B2B9FC2329B6EA7338C3E58705486E95E8E9377B40082;
defparam prom_inst_10.INIT_RAM_30 = 256'hB903CF40DF4DBB7F81D11D27E81C0908C1EB8B0B48C007FF8EA9983F90440ECC;
defparam prom_inst_10.INIT_RAM_31 = 256'h4FE0ABBB9783B624D6EA76F8BDAFF6CC3FC6FA224D4F125E91800FFEAC88B8CA;
defparam prom_inst_10.INIT_RAM_32 = 256'hCCC03FFB7531D6F9D30D10238A72EFE7F7C849D5D35C89A8439E649966201FFD;
defparam prom_inst_10.INIT_RAM_33 = 256'h5DF1ED4B39807FE7F95611A5662EFE2BE3F8DFFC7FB291F4BBD884AF7738E1B4;
defparam prom_inst_10.INIT_RAM_34 = 256'h0ECA058865E75B34E700FFCE6A0C3EBAEEE2DC136328BB288977298677676213;
defparam prom_inst_10.INIT_RAM_35 = 256'h858E1D4F9B1A87A2818EF259CE01FEB8F3D9B1B34EA52FF16D0A72FE633D791C;
defparam prom_inst_10.INIT_RAM_36 = 256'hB06C0FF1737F3AE9DB8368D7D31DC5B39803FD64BB8D85D82B5F3EB0287CE54C;
defparam prom_inst_10.INIT_RAM_37 = 256'hE2D628364CD81864BE1D4F435CC185C22F655E48F83BF605EEFF5BD148279338;
defparam prom_inst_10.INIT_RAM_38 = 256'h8E3A3D91D6C1B47AFA503B4A9D966A1396EEA4867E82BC91E0F7EC0ABC92ABD2;
defparam prom_inst_10.INIT_RAM_39 = 256'h0FDFB0201B320BBDC8FF958CD3206CB322F7D1751762F61F19255363C3EFD804;
defparam prom_inst_10.INIT_RAM_3A = 256'h09CC9B1C7E3F604248285D31C99C4AB040409D8FCCF0A4FDC1D9B90AA6F504C7;
defparam prom_inst_10.INIT_RAM_3B = 256'h53FCC366362B6C78F87EC0AD75FD1329A4F9F14969818C680B8C513350F5105D;
defparam prom_inst_10.INIT_RAM_3C = 256'h03D015B539FFDAA048CDD8F1E0FD806AC8B5F56A6E451B61530216113D7F9874;
defparam prom_inst_10.INIT_RAM_3D = 256'h621F6A39C5761FBAD703ED39B15323E381FB0076B5E0616BF5D9BE6826072684;
defparam prom_inst_10.INIT_RAM_3E = 256'h4D302444F43205FAE4107F4C27D43CC6B1AC67F807F8383CD078BF2706FB5A20;
defparam prom_inst_10.INIT_RAM_3F = 256'h80945B48E084CCA0287F181DB9E7EC22DCD481FD6558CFF00FF0F035DD6B6984;

pROM prom_inst_11 (
    .DO({prom_inst_11_dout_w[30:0],prom_inst_11_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_11.READ_MODE = 1'b0;
defparam prom_inst_11.BIT_WIDTH = 1;
defparam prom_inst_11.RESET_MODE = "SYNC";
defparam prom_inst_11.INIT_RAM_00 = 256'h3FC7C03830745F1611235D5D90D5A90F419E9BB3932BFD1A9AB19FE01FE1E039;
defparam prom_inst_11.INIT_RAM_01 = 256'h964600007E0F80739311FCEB8886BBDFA1CD271FF98B0C9A48D50BE525230000;
defparam prom_inst_11.INIT_RAM_02 = 256'hC3A0122BEC8C0000F03F00666FE4FB9B1EEE774C43A9E3D15B94A3B420B83F14;
defparam prom_inst_11.INIT_RAM_03 = 256'hADF138700891AED79919FE01E0FE01E163E51D878980EE2A87D713AC3F2415F2;
defparam prom_inst_11.INIT_RAM_04 = 256'h1E0EC643ABEE9A6C16E7DD2A3233FC0381F803FD7EA8F1DC0F2DDE310C933587;
defparam prom_inst_11.INIT_RAM_05 = 256'h000000000000055294C8EB9581A82050C71BE00786263BC299E74CA2BE7D668A;
defparam prom_inst_11.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_12 (
    .DO({prom_inst_12_dout_w[30:0],prom_inst_12_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_12.READ_MODE = 1'b0;
defparam prom_inst_12.BIT_WIDTH = 1;
defparam prom_inst_12.RESET_MODE = "SYNC";
defparam prom_inst_12.INIT_RAM_00 = 256'h8FEF0217FFFFFDD607FFFFFF22EFE0000000000000000003F1FFFB0FC7778463;
defparam prom_inst_12.INIT_RAM_01 = 256'hC7FF8C1F9FDF8F0FFFFFF1285FFFFFFE45DF80000000000000000007E3FFE61F;
defparam prom_inst_12.INIT_RAM_02 = 256'h0000003F1FFE180F3FFFED7FFFFFC8F27FFFFF9DBBBF0000000000000000001F;
defparam prom_inst_12.INIT_RAM_03 = 256'h000000000000007E39FC711E3FFF8D5FFFFE0AA47FFFFE3EEF7E000000000000;
defparam prom_inst_12.INIT_RAM_04 = 256'h78F0008000000000000000F8E3F0DA1E3FFF941FFFF860C3FFFFFFFD1CF80000;
defparam prom_inst_12.INIT_RAM_05 = 256'hFFFE0E2BF1E0018000000000000001F1C3E1BC3C7FFF6A1FFFE097C5FFFFFFD5;
defparam prom_inst_12.INIT_RAM_06 = 256'hFE03BD53FFFC005BE3C0030000000000000003E387C27A7CFFFCB43FFF815793;
defparam prom_inst_12.INIT_RAM_07 = 256'hFFF9F2B7BE06CADFFFF807571FE7E60000000000000007C30BC71004FFFA747F;
defparam prom_inst_12.INIT_RAM_08 = 256'h2F1C4003FFEC471F7812EB3FFFF00EAE3FCFCC000000000000000F86178E2009;
defparam prom_inst_12.INIT_RAM_09 = 256'h0000FE185E388001FFECB32EF15FD41FFFE01D5C7F9F98001800000000001F0C;
defparam prom_inst_12.INIT_RAM_0A = 256'h7FFF80000003FC30BC7D40009FAEFB1FE61F203FFFC03B38FF3F30003C3C0000;
defparam prom_inst_12.INIT_RAM_0B = 256'hFCFCC003FFFF0000010FF86178DAC0311F5F6B3FBAFEB07FFFE06671FE7E6000;
defparam prom_inst_12.INIT_RAM_0C = 256'hFFFDABC7F9F9800FFFFE0000063FF0C2F1B580F21F6BCB7F51FF24FFFFF8C4E3;
defparam prom_inst_12.INIT_RAM_0D = 256'hD98617FFFFFF578FF3F3003FFFFC00001CFFE185E36B81E43EF69A7F1DA20FFF;
defparam prom_inst_12.INIT_RAM_0E = 256'h3819D87C0C300FFFF9F8A61FC7038BFFF8F80039FFFF8703C4F7F8601AA2FCFD;
defparam prom_inst_12.INIT_RAM_0F = 256'h13C00000303DEED606F00FFFF7F14C3FCE0703E07FC00071FFFF060789E00000;
defparam prom_inst_12.INIT_RAM_10 = 256'hFFFC185E27803F00202BFD7840601FFFFF86B87FFC07FFE39FFC00E1FFFE0C2F;
defparam prom_inst_12.INIT_RAM_11 = 256'h78000381FFFC38BC4F006300702714B2C4B01FFFFE0D707FF80708383FFC01C1;
defparam prom_inst_12.INIT_RAM_12 = 256'hE0797B04F3C00700FFF873789E008300E0420FF7E9700FFFF81AF07FF07FC77E;
defparam prom_inst_12.INIT_RAM_13 = 256'hC06BC1FFC0FCCC6432E20E01FFF0E6F13C013601E0E70DCAB6F807FFF035E0FF;
defparam prom_inst_12.INIT_RAM_14 = 256'h8FF003FF00D783FF82EC6708DC641C03FFF1CDE27802E403E1879B80FFF003FF;
defparam prom_inst_12.INIT_RAM_15 = 256'h0800AAABC7F801E001AF80FC34F787F3C3E7FE27FFE7E398C8061CDFC3039494;
defparam prom_inst_12.INIT_RAM_16 = 256'hA018FB800003D443AFF001C0035F01F6F60F0FCF0FDCA56FFF8FC031900CD996;
defparam prom_inst_12.INIT_RAM_17 = 256'hF83E018B401217C0002FB2B2DFE031C006BF1FF9933E0F1E3935D59FFE1F00E5;
defparam prom_inst_12.INIT_RAM_18 = 256'h8119AFFFE07847370024D78330DD3775BFC1F300057E3FD249FC0E39C0B91B3F;
defparam prom_inst_12.INIT_RAM_19 = 256'hC7F8311E023FD3FF00F0066600695746619F16687F87E0000BBE001201781C47;
defparam prom_inst_12.INIT_RAM_1A = 256'hA47C7ECE1FF0663905FFAFFE01C00ECC00576F36800C26E0FF1F83E0933C0123;
defparam prom_inst_12.INIT_RAM_1B = 256'hF1FC1383487BF16837E04CE22D097BFC07800D9800859EEC001C0A19FC7E0DC1;
defparam prom_inst_12.INIT_RAM_1C = 256'h181E7CD83C6084DE91FDD3E006AA17E0071E9FE00E003B3465665BBC003A53BF;
defparam prom_inst_12.INIT_RAM_1D = 256'h958F9120383D1CC078C1FDBD23F0BD793FC26FC00E1AFFE01C007668CAC11800;
defparam prom_inst_12.INIT_RAM_1E = 256'h7801D9A3290D3DA01816C440F184FB7A43CF684609D4BF81FC103FE03800ECD1;
defparam prom_inst_12.INIT_RAM_1F = 256'h7844FF80F003B346125526C0382DCDC1C00917F4863DAE9973E97F07FC137FC0;
defparam prom_inst_12.INIT_RAM_20 = 256'hB5A5FC0CF8A7FF01E107668C64911B0071D12083807B2FE90089C2D87FD2FE0E;
defparam prom_inst_12.INIT_RAM_21 = 256'h0FE4DD8CDA89F99C7EBBFE03C20ECD18880714E0011F9C0731215FD203865595;
defparam prom_inst_12.INIT_RAM_22 = 256'hC6ED7F4A19335F01991BF3987CFBFC07841D9A3110115441013A8A0E630CBFA4;
defparam prom_inst_12.INIT_RAM_23 = 256'h0E046E0011F3FEBE1597FF35CC483F540008E007003BE0E56952769B2012201C;
defparam prom_inst_12.INIT_RAM_24 = 256'hBE62B5DAD01140301DE7FD7E5CA1CFF92760FEE80019700E0077C18ADA3C9B85;
defparam prom_inst_12.INIT_RAM_25 = 256'h01DF222B7C4586A0032181FFCBAFFA23655FFFE7DBDFEEF80034201C00EF8115;
defparam prom_inst_12.INIT_RAM_26 = 256'h00FC807003BE4056BC351F036E44C3DE5E5FF471E23FF1BF0CBFDE780067C038;
defparam prom_inst_12.INIT_RAM_27 = 256'h5D1FDC3001F400E0077C80ADFC566196CE99878FABBFE817008E61B8753FBEB0;
defparam prom_inst_12.INIT_RAM_28 = 256'hDFFDE6E7861E9C60038001C00EF9015BFC1F2B2D9C180F13D77FDAD2157FC030;
defparam prom_inst_12.INIT_RAM_29 = 256'hC1FF3E14FCFBCB38E83D3E40057003801DF202B7EC1649001E991E50A4FFBC5B;
defparam prom_inst_12.INIT_RAM_2A = 256'h39565C0E31FD4889FFFF82DB50A8D2C87EC91F80337005CFF8186A601EEA39EB;
defparam prom_inst_12.INIT_RAM_2B = 256'hF0FF088018FD8FB193FD94C3FFFF0A67F40611F07DB42F0066E00B9FF4731750;
defparam prom_inst_12.INIT_RAM_2C = 256'hBB802E7FE1EA810001CEF1CF27E99BE7FFE0032C707B60E0FB165E00DDC0173F;
defparam prom_inst_12.INIT_RAM_2D = 256'hA4CFF00373005CFFFC2DA2403A84B61E4FDF405FFFC022127DA58101F5E4B801;
defparam prom_inst_12.INIT_RAM_2E = 256'hE7C1E1036A73E006E600B9FFF80E940075506B021FACEE7FFC0008F896920203;
defparam prom_inst_12.INIT_RAM_2F = 256'hC01ECA0893A1F806C847800DCC0173FFF028A0000EBFB51C3F1102FFF00098E7;
defparam prom_inst_12.INIT_RAM_30 = 256'hFFF3F7FF803F681F067CFC0EA81F001B9802E7FFE1EA43011EF3793A7E3A13FF;
defparam prom_inst_12.INIT_RAM_31 = 256'h7C46B6E8F207FA20D343886A34342A0B66CF083B28C5D01FC2E50780AA2CF8C8;
defparam prom_inst_12.INIT_RAM_32 = 256'hFC5E8030C0F42969DC3FF331498B100EBE816E36F9DE1076D18BA00FFE2A51D5;
defparam prom_inst_12.INIT_RAM_33 = 256'h4F2E003FF89D2C9086EC0661F19FF3F06F89D6CF5493CC2CAE3C20EDA717001F;
defparam prom_inst_12.INIT_RAM_34 = 256'h8F7001B6BE5C007FF1AB0BA04C7E240027FFF9A277B6F5E9909F8059807800DB;
defparam prom_inst_12.INIT_RAM_35 = 256'hAA1F69E1EEC003697CF800FFF39AC74118FFDB162880435BB8E419B5961BB7B3;
defparam prom_inst_12.INIT_RAM_36 = 256'h01134DF16CB231D1CF8006D3F9F001FFFF140F0379F001306F0036C235139466;
defparam prom_inst_12.INIT_RAM_37 = 256'h2C0052D2071124B1EFDBF93D93000DA7FBE003FFF11F0701D7FCF693D8010484;
defparam prom_inst_12.INIT_RAM_38 = 256'hB9FFC2CA773E7782F999B971ED35F7F818003B4FFBC007FFE33F1513BF9FC4CF;
defparam prom_inst_12.INIT_RAM_39 = 256'h0A1518F96DFFC372E2EFEE00E8EF0D13A329A3003000769FF7800FFF8722757C;
defparam prom_inst_12.INIT_RAM_3A = 256'h9E003FFE1516B0E1A6BFD14A94FBE007DFEB52E60C7947426000ED3FCF001FFF;
defparam prom_inst_12.INIT_RAM_3B = 256'h0001B4FF3C007FFC234261DAE03FE98D3623802B17ADE6CC654BEA808001DA7F;
defparam prom_inst_12.INIT_RAM_3C = 256'h8AABB270000369FE7800FFF80A84185B0B7FEE1F931207FAB8D95FC93F3CC929;
defparam prom_inst_12.INIT_RAM_3D = 256'h5BC9C902CFD0AAC00006D3FCF001FFF06848707B45FF03EFA6F00C03203A9F53;
defparam prom_inst_12.INIT_RAM_3E = 256'h41EBFC3000C8DAF57AE26480000DA7F1E003FFE0C8E2E174F7FF189167FC7EED;
defparam prom_inst_12.INIT_RAM_3F = 256'h3F7F071AFC68DECB4A71E33B0DF5CFC0003B43F5AFFFFFC1F6B558566FFC1C53;

pROM prom_inst_13 (
    .DO({prom_inst_13_dout_w[30:0],prom_inst_13_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_13.READ_MODE = 1'b0;
defparam prom_inst_13.BIT_WIDTH = 1;
defparam prom_inst_13.RESET_MODE = "SYNC";
defparam prom_inst_13.INIT_RAM_00 = 256'hF0968E458FFF0F003B2921CDDC04F3FAE49BE7A0007687EB500FFFFFFBED9303;
defparam prom_inst_13.INIT_RAM_01 = 256'h003FFFFFEB5D8B2DBC5E1FF4A98AF6DCE290218850A3364000ED0FDC801FFFFF;
defparam prom_inst_13.INIT_RAM_02 = 256'h03B47FB2007FFFFFD5802B5751BE03C16AFCF2E45477C1AC6230EDC001DA3FF9;
defparam prom_inst_13.INIT_RAM_03 = 256'h39C456000768FF4400FFFFFF86031E44457E71D73F4237789929602D5FE32A80;
defparam prom_inst_13.INIT_RAM_04 = 256'h5B68062EF156EC000ED1FE8801FFFFFFD61636D9EEFEF0912E32F060EA99C788;
defparam prom_inst_13.INIT_RAM_05 = 256'h0562008F272707F2DD608C001DA3FD1003FFFFFEAA0CB84177FF801F38390AB4;
defparam prom_inst_13.INIT_RAM_06 = 256'hD78B860604D036BC151B0ADF037A40003F57FA5007FFFC03DF2C20A7F3FC0003;
defparam prom_inst_13.INIT_RAM_07 = 256'h16B0FF4A3A7EBE007E0DC8193536BE7B6DD4E0007EAFF4E00FFFFF0529807C38;
defparam prom_inst_13.INIT_RAM_08 = 256'hFFFFF8028680FBA0FFFF7FE9F7682859F4180ECE8508C000FD5FE9C03FFFFC02;
defparam prom_inst_13.INIT_RAM_09 = 256'hBD7FB303FFFFE003CDC02FA63F0C1FF93D522DD1A2FB5E2FE28CC001DABFD380;
defparam prom_inst_13.INIT_RAM_0A = 256'hF0A300077AFFE60F7FFF8007D20007B1C9303FFB8BD3590BC8D88B2499A88003;
defparam prom_inst_13.INIT_RAM_0B = 256'h0943317BEA94000EF5FFC83EFFFF00085F80731DBC953851FB044CF73A0E937F;
defparam prom_inst_13.INIT_RAM_0C = 256'h782656329121D4487820001DEBFF907DFFFE008A7182A8CD8E6A7132640B4AE2;
defparam prom_inst_13.INIT_RAM_0D = 256'hBBB9C002426446E9335F8054D2380860B7FBC8FBFFFC014CA30C6278FE00E292;
defparam prom_inst_13.INIT_RAM_0E = 256'h6770F240783F8D960F58E56AA146A230477000C16FF791FFFFF807CDC3B87BA1;
defparam prom_inst_13.INIT_RAM_0F = 256'hFF8001E266E0EFEAE403FB321B9C7AFCACA9317D56E00182DFEF03FFFFE001A4;
defparam prom_inst_13.INIT_RAM_10 = 256'h7FFA0FFFFE0003594C60EE0720FF0E27EA3C63DD5A77D1985FC00305BFDE07FF;
defparam prom_inst_13.INIT_RAM_11 = 256'hC7000C16FFA61FFFF000063B0460EB55D21C1E3C407D9D04940888909380060B;
defparam prom_inst_13.INIT_RAM_12 = 256'h2BF4D66F8800182DFF4C3FFFC0000CEB0CE09BCB988CE0E03F57DC13247CB91B;
defparam prom_inst_13.INIT_RAM_13 = 256'h83907A4FDA87C7F51000305BFE987FFF0001095C19E1C8F45387F18CB712FF66;
defparam prom_inst_13.INIT_RAM_14 = 256'h37831637D5BA07740B1E3E1A140030B7F7307FFC000203EC3BC31CC5B4009761;
defparam prom_inst_13.INIT_RAM_15 = 256'h45824FEBBF0535E6586EF1E6F762DCCC4800656FEE60F7FF870409C8C6C136DB;
defparam prom_inst_13.INIT_RAM_16 = 256'h001FF9C4CF0413E01F0D08B107CAF95D6E1286107800CEDFD4C0EFFF0000FD9B;
defparam prom_inst_13.INIT_RAM_17 = 256'h5303BFE003C039229E4874B53E0B47C2444C54E79F6BEE4130419DBFA981DFFC;
defparam prom_inst_13.INIT_RAM_18 = 256'hC1077EEFA6037FFF7C000815BDC2C318FC1AA797CBD6EA72489D5F82E083BF7F;
defparam prom_inst_13.INIT_RAM_19 = 256'h46D34F81820EFDDF4E06FFFF001F0AB13F8B5A51F83472F85C95B685819B4E81;
defparam prom_inst_13.INIT_RAM_1A = 256'h779D0C555ADB047F0C1DFB9E9C0DFFE001F1662B7F1FFF43F84F7A81BF58880B;
defparam prom_inst_13.INIT_RAM_1B = 256'h831B36B65D93A4A6021D6DD71833B43C3003FF003F82C6BEFE2CC317F1833F62;
defparam prom_inst_13.INIT_RAM_1C = 256'h3516D50F067F3A282715A8F383ADAFAE3067687860070784700586489AB569DF;
defparam prom_inst_13.INIT_RAM_1D = 256'h0004C9A37E21C17C0DD4BDE8B961FBCFB441A75C20CED0F0C0100E01C0002FD1;
defparam prom_inst_13.INIT_RAM_1E = 256'h003FC03C00DC05C2EAC8A7403379F7161E1C685514CF8230419DA1E180200007;
defparam prom_inst_13.INIT_RAM_1F = 256'h0672878600FF83F81FB9BE8799A961800082EFB61674F7E40BC44C60833B43C3;
defparam prom_inst_13.INIT_RAM_20 = 256'h215723800CE50F1C00FC3FFEFF72682F3BF98DF832A7BCA002FAB738F4A6B0C0;
defparam prom_inst_13.INIT_RAM_21 = 256'h2E7DA9B0AD33030019CA1E3801F1FFFFFFC66C4E003EB9F89077C98BED0EE192;
defparam prom_inst_13.INIT_RAM_22 = 256'h702839F3BDC6DFD81F18B3F81BF63CD07BC3FFFFFF18A8DCA89BF7FB97161B02;
defparam prom_inst_13.INIT_RAM_23 = 256'h96CDA9F33A0AFD954A1E8EDB59FD572077E879A0333FFFFFFFE590D483519BCD;
defparam prom_inst_13.INIT_RAM_24 = 256'hFFC72154ECFD618107A8F3790CDD4AF05FF6A220CFD0F2981F8FFFFFFFCF91A8;
defparam prom_inst_13.INIT_RAM_25 = 256'h3F000FFFFFEC827E90BF850208CCE2A81261112F525C35819FA1E57C3FFF1FFF;
defparam prom_inst_13.INIT_RAM_26 = 256'h7E0797F003000FFFFFFBC0EEBCF87C41C8261A3A804D9562AB49A4833F03CAFC;
defparam prom_inst_13.INIT_RAM_27 = 256'h078494E6FC0725C139E00FFFFF5481BCA9E96B0850A5B698370E282A4E129103;
defparam prom_inst_13.INIT_RAM_28 = 256'h431B4937CED4EFE5F80E6A0059E00FFFFEBB0325427FBF2918AC917E0290FB33;
defparam prom_inst_13.INIT_RAM_29 = 256'h566DBCCBD873E0591E732264783C4F0A43C00FFFFE42022187BB65423E446346;
defparam prom_inst_13.INIT_RAM_2A = 256'hCD743678E02C80A9F82DADE0EA3B3288F0789E3893F43FF8784347D6E673EB3F;
defparam prom_inst_13.INIT_RAM_2B = 256'hFC108989F9DC54DC2599980583310034498DA531E0F57C7CACEC3FF0F4D10D65;
defparam prom_inst_13.INIT_RAM_2C = 256'hC43801C3F8294553D02CA8341D8CF9DC766FD57F98D65A63C1EAB8FE70F823E1;
defparam prom_inst_13.INIT_RAM_2D = 256'h07B538FE7C780007D4CA15A770FBA074A67CEE4721EB16A163D49FC783D2784F;
defparam prom_inst_13.INIT_RAM_2E = 256'h635FD31E0F6A1FFC0CF8000FF155B2EE134641EFA03D425347FEF395768DBF8F;
defparam prom_inst_13.INIT_RAM_2F = 256'h5EEAEE88BFAABE3C1ED71FF80078001FFB679D5F0F2CA2AD1D7A0081CD3A010D;
defparam prom_inst_13.INIT_RAM_30 = 256'h3CDD43A87DB7C3E003E613081D983DE44CF8003FC62F3AF578564F2C62F42F42;
defparam prom_inst_13.INIT_RAM_31 = 256'h21702368313A30C15AEA5D125A0F96103B3011C029F8007A56F032D7D0B011A6;
defparam prom_inst_13.INIT_RAM_32 = 256'h975FCF78A3E052C06274CDF2ABE5F31AE71DAC20F67E018044F000F66FCA45AC;
defparam prom_inst_13.INIT_RAM_33 = 256'h2F2001F43E251C93631474C0CDCD78DF754E1A49A6DC5841EEBF3800EAC001FE;
defparam prom_inst_13.INIT_RAM_34 = 256'hFA3FFC00057001E9FE6B18A6E6FCEDC39312BCEA4E755ABE15BE31837D1FF800;
defparam prom_inst_13.INIT_RAM_35 = 256'hF868C51DB4FDFE0052F003F28F0014ADC6FDE9FE64259FC9E00A807B64526306;
defparam prom_inst_13.INIT_RAM_36 = 256'h61E62CC62C39AA316BF38710B3F003E74B5C2F598FFAD2F9D854E0A462FDD173;
defparam prom_inst_13.INIT_RAM_37 = 256'h6333D5070C790E53C69510FEA8E70F20B7E003BE97AA5D9B1FF5B063B2E9B593;
defparam prom_inst_13.INIT_RAM_38 = 256'hE78440F8C66DEA81120AD52F29AC21FC53CFF924AF003BFE7D298224E71A187C;
defparam prom_inst_13.INIT_RAM_39 = 256'h1E265C8054C443E18DC1459D67A3B9CFBD7443F9A79FF2018E0073F432732A4B;
defparam prom_inst_13.INIT_RAM_3A = 256'h98004FFA1C34FC89EB088FC73B9F089A97A68E00F59E47F3CE3FE400CC0067EA;
defparam prom_inst_13.INIT_RAM_3B = 256'h78FFFE5E30000FFA41E8B15C7C81BF0C769CD58569EDB81A65540FE39C7FDC22;
defparam prom_inst_13.INIT_RAM_3C = 256'h4E7C3F86F1FFFEB160001F2CCAD9B33A6233FC18EDCC693FBC85B01E25681FFB;
defparam prom_inst_13.INIT_RAM_3D = 256'h4697B3A4B9807E7DE2018EC8E0003E4CB5F7DA37B0ABF031D2325F76C844411E;
defparam prom_inst_13.INIT_RAM_3E = 256'h01CA71A8FB346CC713A9E366F4031D99C0007DC6DBED70285957E0E3A07FA700;
defparam prom_inst_13.INIT_RAM_3F = 256'h10FF070E031F6E71CC34FD9E3751C6CFE00006936000FB2A03A3018A5C7FC3C3;

pROM prom_inst_14 (
    .DO({prom_inst_14_dout_w[30:0],prom_inst_14_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_14.READ_MODE = 1'b0;
defparam prom_inst_14.BIT_WIDTH = 1;
defparam prom_inst_14.RESET_MODE = "SYNC";
defparam prom_inst_14.INIT_RAM_00 = 256'hD5D2F642E3DE0E164EA7425C25AD3E354EA39EAFC0000D2CC001FE7F36C00A92;
defparam prom_inst_14.INIT_RAM_01 = 256'h0003F088ED27E76CCFF07C0CED2E84688446D5079D472D5EC0001A718003FCD3;
defparam prom_inst_14.INIT_RAM_02 = 256'h0000710E0007F025D81CE2721F83F811DD60363E88AD29D3BA8F5A99800038C7;
defparam prom_inst_14.INIT_RAM_03 = 256'hEA3ED8020000929D000FE61790226B8B000FF023FF760FEE210CBF6E751EF531;
defparam prom_inst_14.INIT_RAM_04 = 256'hE32224F1D47DB2040001257A000EEEDF088ACD9A003FE01E7F916EC9C465ECD4;
defparam prom_inst_14.INIT_RAM_05 = 256'h0D1D94FBE400BF9F107B7078000244B4001DD55A81ABFAC43C7FC57C8CB722BC;
defparam prom_inst_14.INIT_RAM_06 = 256'hE46E35CA1BBB169CA6DB76A4E0F6B1F00001E94800071E825576A4BF1FA78AE1;
defparam prom_inst_14.INIT_RAM_07 = 256'h003ED4E1C79CF9D4ADF71C82D559E44241EB67E00003D290001E300AD0EC596F;
defparam prom_inst_14.INIT_RAM_08 = 256'h00FC3C67AD712B8E3421E8A77B44649AC79DD72B43D53FC02004AD20007E2677;
defparam prom_inst_14.INIT_RAM_09 = 256'h0001728003F80595DE5BA447CC07588FD4521F65AADF08DC03AA7F81C000BB40;
defparam prom_inst_14.INIT_RAM_0A = 256'h0F59F100000125000FFE45BCB5603CC0BD1C750F9CA3231ED290E4DF0774FC00;
defparam prom_inst_14.INIT_RAM_0B = 256'hA11FA7801EA3C3F8001A4A001FFEA8034B05F4385E70B85E98F8E1CCEE7E5972;
defparam prom_inst_14.INIT_RAM_0C = 256'h797FC7420EB71528117007FC003494003FFD60A607F4F0F35CE13ABD7AB693FE;
defparam prom_inst_14.INIT_RAM_0D = 256'hC43FA7F0FD46F5A215F2EA5022A007E00660BE1FFFC3974D8C75BF87F20AC3F8;
defparam prom_inst_14.INIT_RAM_0E = 256'h322FF99F18BDAFE1F89CE567178E74A0442000000CC57C1FFF872F9B1F18C00F;
defparam prom_inst_14.INIT_RAM_0F = 256'hFE3B0F8E03B684FC31AFDF03E77CF893A31369409D80000011DA783FFF1E8736;
defparam prom_inst_14.INIT_RAM_10 = 256'h479DF0007C75DF1E2FF9077824F13C07EC3C3B15CD9652813F8038002384F83F;
defparam prom_inst_14.INIT_RAM_11 = 256'hB20183000FFBE000F8FF280D065F0771A9AFF90F401BF0B4D777A50259008000;
defparam prom_inst_14.INIT_RAM_12 = 256'hE11A949B58023E001EF3C001F1EE518A4EBC1EE79385E61F7C2E57019B0F4A44;
defparam prom_inst_14.INIT_RAM_13 = 256'h0AB6E9724C2A2995F4E558003DF78003E1DCAB153C4F30CC6BAFCC3CA34CAA26;
defparam prom_inst_14.INIT_RAM_14 = 256'h5BFD906F2B50A4A72AEAF3E84FCB26403A578000943D25D5E6F8BF310DFEC831;
defparam prom_inst_14.INIT_RAM_15 = 256'hC36663FAE7F321D3A9BC7FB8851487C4270CE210729F003ED8784B68A9713CB7;
defparam prom_inst_14.INIT_RAM_16 = 256'h49E12406341C0FC95FE003E2469ACF58E2501FBBD80150A0212E2FDE52F0924D;
defparam prom_inst_14.INIT_RAM_17 = 256'h480060182B43C9C84A7073B56F8005F034A94D6661A43F7626218240340F01C2;
defparam prom_inst_14.INIT_RAM_18 = 256'h7517F8079DF0FF8FD687C5B45400E0171E0002E2CA962C44EEB87E1CCCB66600;
defparam prom_inst_14.INIT_RAM_19 = 256'h2F85F1977433AC1E1C7EF0E99D0E417AD9FFC7EE340004AFF7DB8818DC88F8D0;
defparam prom_inst_14.INIT_RAM_1A = 256'hA6D2A373DF77EBC8467A007F4400C42FBA1F38AB9FFE31D068001886EB7A59BC;
defparam prom_inst_14.INIT_RAM_1B = 256'h2185ECB72ECE8C458FDFD784777AD8AC30C8C3F47802F78F4BF71B2080D03927;
defparam prom_inst_14.INIT_RAM_1C = 256'h27FC3F62031BC723C76724F9ECCFA96DEE7B115313231F88D46D2E3C93FE3EB2;
defparam prom_inst_14.INIT_RAM_1D = 256'h73FB71E647FC3B088201DB89DD3CEA53F61F233B2F36460159BCFC111EB07CF9;
defparam prom_inst_14.INIT_RAM_1E = 256'h870F01F8CE68078CCFF872310003A9B775409B135A3A454A49185C150C43E075;
defparam prom_inst_14.INIT_RAM_1F = 256'hEDC8742E567F810046A61C31CFF0FF6820DA0F83B4A07CB7FC3606B655116810;
defparam prom_inst_14.INIT_RAM_20 = 256'hA48969A4B5F37810A1FFC163A31C70E39FF18E2441F48E78843DF34B50448BE8;
defparam prom_inst_14.INIT_RAM_21 = 256'hCA33BCDB7913ED6566777171C3FFC2E49ACCE3C73FE119C8801C6E5E514EACC8;
defparam prom_inst_14.INIT_RAM_22 = 256'hB90FC54147220AC48227D8C8DA8A5829EFFE021DC8E39F183FE58DF15F6FF52E;
defparam prom_inst_14.INIT_RAM_23 = 256'hFF823EE3428D9319F39BFFA8044FF921E5F3910BDFFC04BB11C73E307FC918B2;
defparam prom_inst_14.INIT_RAM_24 = 256'hC738F1C3FF04DAC6383558AD90BDDD58408BB1438CE1FBD3AFF81BAA038E78E0;
defparam prom_inst_14.INIT_RAM_25 = 256'h0FE07B0D0E738787FE01968C525FD828304C406101077903FC7331BD0FF02F90;
defparam prom_inst_14.INIT_RAM_26 = 256'h6DF07AED0FC0296A18E70E0FFCC5121998BC7A89DC82BCCC020E82837CDE724F;
defparam prom_inst_14.INIT_RAM_27 = 256'h085ECC3C4B5CFCCA1F80DAA031CE381FF9CB6E12E2B37A708768C936040F7902;
defparam prom_inst_14.INIT_RAM_28 = 256'h5AFFE6E917B72C529BD7D3D41F02A324639C707FF3D65425451DD23D7854235C;
defparam prom_inst_14.INIT_RAM_29 = 256'hC0DB29FD3637F03227EE960E6C5BFED87FFF0551C670E3FFFE7C61F6413D5F92;
defparam prom_inst_14.INIT_RAM_2A = 256'hF9CBF0C8B2C79A6AEDE0F5844FD72C0E9501AC30FFE9A2A38CC3CFFFFCF2C7EF;
defparam prom_inst_14.INIT_RAM_2B = 256'h230E3FFFD25A99213FACD36C8F30CBC89EA45C0E48934441FF9E44C719879FFF;
defparam prom_inst_14.INIT_RAM_2C = 256'hFC0CCCB88C3C7FFFB625C03819B2BBD7F9700D9120C098D2805657C3FE0EAD4C;
defparam prom_inst_14.INIT_RAM_2D = 256'h1B88081FF039F9F118F0FEFFE7AA70BD17FF63E979388C2241BCF9AB18AC6F87;
defparam prom_inst_14.INIT_RAM_2E = 256'h7752F0985A12C43FE05915E631E1FDFF8508E8BB8E58B1A35CB930458B79F92A;
defparam prom_inst_14.INIT_RAM_2F = 256'hF01BE1285B94F123BC25BC7FC3D32F8CC7C3F3FF099252153B48C2581A4FBC8B;
defparam prom_inst_14.INIT_RAM_30 = 256'h8F49B0C7D81D7354D629FFF2C4E8EE88FC1C0A138F07FFFFD1525801912D6C27;
defparam prom_inst_14.INIT_RAM_31 = 256'h71303822A6F6F02B305AC6AAA85FF0577620CD3378F0146F1E0FFFFF36D7B808;
defparam prom_inst_14.INIT_RAM_32 = 256'hF0FFFFFC556F70CB4D2EB215C871CF5654246A5692E06FD296E068DE783FFFFE;
defparam prom_inst_14.INIT_RAM_33 = 256'hD981CE73C1FFFFF8157171A02B647CDBF5231E933058D794C50DE8CA6440F138;
defparam prom_inst_14.INIT_RAM_34 = 256'h0F90697801079DC707FFFFF108DDFE2C97C074A68A973D3A24C1E662C32DAB63;
defparam prom_inst_14.INIT_RAM_35 = 256'h72E1F04BC570466FDA0F7B9E0FFFFEC62805C9AF480E1FB4A06C7AE538B1F5B7;
defparam prom_inst_14.INIT_RAM_36 = 256'hC48021E8F9A27225B22563B27C1EF63C1FFFFD9CEC3913AF3DB0FF3EC4F4F5FA;
defparam prom_inst_14.INIT_RAM_37 = 256'hC2544D341080445E82F627D3077654BC50799870FFFBFFF93C0EE5707AB2BABC;
defparam prom_inst_14.INIT_RAM_38 = 256'h9C1B1F916F17147A42408C2B973429EE4541D27900F330E1FFF7FFFCE7FE2EFE;
defparam prom_inst_14.INIT_RAM_39 = 256'hFFDFFFE3D00A766924C1BC8AC1810E4FD583B83C125F4DEEA1C66383FFEFFFF9;
defparam prom_inst_14.INIT_RAM_3A = 256'h8E771C1FFE3FFFCCCE6B2FCE8B7A7B955102046A832B9E7C6B8577DBC739C707;
defparam prom_inst_14.INIT_RAM_3B = 256'hB1033CFB38CC707FF87FFF50CDA0DEFDB1AD7397D204BCAF4EA79E9CAE0C8FDF;
defparam prom_inst_14.INIT_RAM_3C = 256'h19F57D92FDFE23A27111E0FFE0FFFFBC9F3BE87743AD07BCDC097EBBA454F576;
defparam prom_inst_14.INIT_RAM_3D = 256'hD4365F1E434F00AE7B000FF5C263C3FF81FFFC05675AD50D8DCC041DD811FE22;
defparam prom_inst_14.INIT_RAM_3E = 256'h0F478E1EF86C69BED95CF2A5F7E7D63F3ECF87F807FFC039A2F98D88B3C02F08;
defparam prom_inst_14.INIT_RAM_3F = 256'h15B7A3ED3CAA7C34B0C62D4582815B409CE7284E799F0FF00FFF003695B01091;

pROM prom_inst_15 (
    .DO({prom_inst_15_dout_w[30:0],prom_inst_15_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_15.READ_MODE = 1'b0;
defparam prom_inst_15.BIT_WIDTH = 1;
defparam prom_inst_15.RESET_MODE = "SYNC";
defparam prom_inst_15.INIT_RAM_00 = 256'h3FF8003FDBDBC070F9FC784061AD9D876697EB1E902CA01CE33E1FE01FFE003E;
defparam prom_inst_15.INIT_RAM_01 = 256'h187800007FF0007C18A6A1A88622F09FC37EC40F769C0911071970F9C63C0000;
defparam prom_inst_15.INIT_RAM_02 = 256'h3CC593CCF0F00000FFC0007876A67226A750E10786D3383F169A66DA9F22A9E7;
defparam prom_inst_15.INIT_RAM_03 = 256'hCF3178E1F11BAF19E1E00001FF0001FE7752E84EB7C7C38D0D41E033D67C441E;
defparam prom_inst_15.INIT_RAM_04 = 256'h36B09E003DA278D3E4F4DE33C3C00003FE0003FE6B81DCE3F48F84C21A91D2A1;
defparam prom_inst_15.INIT_RAM_05 = 256'h00000000000008D8743D5CDC2DF8386707E00007F9C03BFCD83F6F10E8E642C4;
defparam prom_inst_15.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_16 (
    .DO({prom_inst_16_dout_w[30:0],prom_inst_16_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_16.READ_MODE = 1'b0;
defparam prom_inst_16.BIT_WIDTH = 1;
defparam prom_inst_16.RESET_MODE = "SYNC";
defparam prom_inst_16.INIT_RAM_00 = 256'h0FEF0EF7FFFFFE37FFFFFFFF3B1FE0000000000000000003FE00035807F7842A;
defparam prom_inst_16.INIT_RAM_01 = 256'hF8000D601FDF99FFFFFFFE6FBFFFFFFE763F80000000000000000007FC0006B0;
defparam prom_inst_16.INIT_RAM_02 = 256'h0000003FE0001AC03FFFE1FFFFFFFC9F3FFFFFFDDC7F0000000000000000001F;
defparam prom_inst_16.INIT_RAM_03 = 256'h000000000000007FC00074803FFFF51FFFFFF1FF7FFFFFFF30FE000000000000;
defparam prom_inst_16.INIT_RAM_04 = 256'h87F0008000000000000000FF0000F1003FFF241FFFFF83F9FFFFFFFE63F80000;
defparam prom_inst_16.INIT_RAM_05 = 256'hFFFE0E320FE0018000000000000001FE0001EA007FFE801FFFFF13EFFFFFFFD9;
defparam prom_inst_16.INIT_RAM_06 = 256'hFFFC9FAFFFFC006C1FC0030000000000000003FC0003D600FFFF043FFFFE3FFF;
defparam prom_inst_16.INIT_RAM_07 = 256'hFFF61A37FFF97DBFFFF80798FFE7E60000000000000007FC00074800FFFD947F;
defparam prom_inst_16.INIT_RAM_08 = 256'h001D2003FFF3A41FFFE1F1FFFFF00F31FFCFCC000000000000000FF8000E9001;
defparam prom_inst_16.INIT_RAM_09 = 256'h0000FFE0003A4001FFF3702FFF8BEFFFFFE01E63FF9F98001800000000001FF0;
defparam prom_inst_16.INIT_RAM_0A = 256'h7FFF80000003FFC00078C0009FF0581FFF1FEFFFFFC03DC7FF3F30003C3C0000;
defparam prom_inst_16.INIT_RAM_0B = 256'hFCFCC003FFFF0000010FFF8000F1C0011FE0983FBC1F6FFFFFE07B8FFE7E6000;
defparam prom_inst_16.INIT_RAM_0C = 256'hFFFDCC3FF9F9800FFFFE0000063FFF0001E380021F9C197F7A7D5FFFFFF8F71F;
defparam prom_inst_16.INIT_RAM_0D = 256'h0F35F7FFFFFF987FF3F3003FFFFC00001CFFFE0003C780043F391E7FE3B9FFFF;
defparam prom_inst_16.INIT_RAM_0E = 256'h37FE387F0CC7FFFFF9FF39FFC70383FFFFF80039FFFFF80007AFF8001F7F1CFE;
defparam prom_inst_16.INIT_RAM_0F = 256'h1EA000002FFE1CE8A76FFFFFF7FE73FFCE0F03EFFFC00071FFFFF8000F500000;
defparam prom_inst_16.INIT_RAM_10 = 256'hFFFFE0003D403F001FEC1D814E1FFFFFFFF8C7FFFC07FFFF9FFC00E1FFFFF000;
defparam prom_inst_16.INIT_RAM_11 = 256'h00000381FFFFC0007A807F000FF8FD45DB4FFFFFFFF18FFFF8070FF83FFC01C1;
defparam prom_inst_16.INIT_RAM_12 = 256'hE0FED7F8FC000700FFFF8000F500FF001FFDDF8BFA8FFFFFFFE30FFFF07FFD00;
defparam prom_inst_16.INIT_RAM_13 = 256'hFF8C3FFFC0FC49F83D020E01FFFF0001EA01CE001FF89D1AC907FFFFFFC61FFF;
defparam prom_inst_16.INIT_RAM_14 = 256'h400FFFFFFF187FFF833478F0E3841C03FFFE0003D4031C001FF81EA1600FFFFF;
defparam prom_inst_16.INIT_RAM_15 = 256'hF7FF0F0C0807FFFFFE307FFC3F3FF803FC07FDB7FFF8001F980704183CFC1716;
defparam prom_inst_16.INIT_RAM_16 = 256'hE01D581FFFFC3C50100FFFFFFC60FFF7F70FF00FF013356FFFF0003F300EC819;
defparam prom_inst_16.INIT_RAM_17 = 256'hFFC001F5C018B03FFFF032C9201FCFFFF8C0FFFFE01FF01FC033E59FFFE000FA;
defparam prom_inst_16.INIT_RAM_18 = 256'h019FEFFFFF8047CA8032B07CCFE247E2403E0FFFF981FFFD01FFF03E00F8C33F;
defparam prom_inst_16.INIT_RAM_19 = 256'hC7FFC1E003FF13FFFF000795004630B99FE0370780781FFFF201FFE201FFE078;
defparam prom_inst_16.INIT_RAM_1A = 256'hC803804A1FFF87C007FE2FFFFE000F2A008B21797FF3B71F00E07C1FE403FEBC;
defparam prom_inst_16.INIT_RAM_1B = 256'h0E03E07F9004038807FF8F000DFA5BFFF8000E5401334273FFE331E60381F03F;
defparam prom_inst_16.INIT_RAM_1C = 256'hE7E1DF37C39F05FF2003370006DC180007E11FFFF0003CAC063CC6A3FFC177C0;
defparam prom_inst_16.INIT_RAM_1D = 256'h18FA9C3FC7C2DF3F873EFBFE400A47E83FFC70000FE53FFFE00079580C7A8897;
defparam prom_inst_16.INIT_RAM_1E = 256'h8001E56033F9093FE7E867BF0E7917FC8009CF5E0FF8C001FFEBBFFFC000F2B0;
defparam prom_inst_16.INIT_RAM_1F = 256'hFFCAFFFF0003CAC027F7287FC7D1AB3E3FF50FF90027F75F1FF18007FFE47FFF;
defparam prom_inst_16.INIT_RAM_20 = 256'h76C6000FFF9BFFFE000795804FFB767F8FA06F7C7F951FF20081FDEFFFE3000F;
defparam prom_inst_16.INIT_RAM_21 = 256'h0E2F26713D0E001FFF45FFFC000F2B00DFEBFDFFFFE013F8CE123FE403B43AE6;
defparam prom_inst_16.INIT_RAM_22 = 256'h3BDCFF921CB6E0FCBE1C001FFF83FFF8001E5601BFE6FA7FFFC5D7F19D9E7FC8;
defparam prom_inst_16.INIT_RAM_23 = 256'h9FF879FFE439FF28EC8800C15B77C077FFF2AFF8003CA80639A548E7DDCCBFE3;
defparam prom_inst_16.INIT_RAM_24 = 256'hFFCDE9E73FE2FFCFD473FE5F8DDE0006B99F00EFFFE5FFF00079500C7BDBC8FB;
defparam prom_inst_16.INIT_RAM_25 = 256'h01E56031FFCBDEDFFFC1FE0064E7FCBDF7A00018A6C000FFFFCCFFE000F2A018;
defparam prom_inst_16.INIT_RAM_26 = 256'hFF09FF8003CAC063FF9BC7FF9F82FC20B1CFF95A3FC0006C7940007FFF9D7FC0;
defparam prom_inst_16.INIT_RAM_27 = 256'h2A00003FFE01FF00079580C7FF19A7EF3F45F872879FF2FD7F7000006E8000BF;
defparam prom_inst_16.INIT_RAM_28 = 256'h800206E0E401007FFC1FFE000F2B018FFE10FFDE7FA9F0E68F3FEF79E2800000;
defparam prom_inst_16.INIT_RAM_29 = 256'h24FFA89733000F396402007FF857FC001E56031FEC19BFFFFF65E193167FD6FF;
defparam prom_inst_16.INIT_RAM_2A = 256'hFA8F1D59FBFC73BE000003DF67D40CFF806AA0003CA806BFF813839FFD27C258;
defparam prom_inst_16.INIT_RAM_2B = 256'hF0F1F7FFFF0173C617FEBCFC000003EFF50801FF80B3D00079500D7FF07953EF;
defparam prom_inst_16.INIT_RAM_2C = 256'hC54035FFE1F173FFFE0B1FD02FFDCFD8000003EFE3E300FF01C4A000E2A01AFF;
defparam prom_inst_16.INIT_RAM_2D = 256'h020200038A806BFFFC3347BFDD112CC05FFE27A0000023DDD26401FE00094001;
defparam prom_inst_16.INIT_RAM_2E = 256'h1E41E1FC062C00071500D7FFF8132FFFBA607452BFFD318000000F87E64083FC;
defparam prom_inst_16.INIT_RAM_2F = 256'h001FCDF06861F9F80578000E2A01AFFFF037FFFFF0DFB4377FED390000009F18;
defparam prom_inst_16.INIT_RAM_30 = 256'hFF730800003FEFE17BF8FFF02360001C54035FFFE1F7BEFFE17FC42CFFC26400;
defparam prom_inst_16.INIT_RAM_31 = 256'h8009DF4DF7D001C4107FFFF40344EBC05A10003CB806901FC3FCFC7D45C7C079;
defparam prom_inst_16.INIT_RAM_32 = 256'hFC6C9FCF0003C79259E0030051F7FFF88541FFC080200079700D200FFE328E23;
defparam prom_inst_16.INIT_RAM_33 = 256'hC034003FF8EC1F7F0703E8DBF5C012400FF7EF3C9753FFC021C000F2E01A001F;
defparam prom_inst_16.INIT_RAM_34 = 256'h680001CB8068007FF1DD3C7F6F81D385BE0022407FE28E17B37FFF80DB8000E5;
defparam prom_inst_16.INIT_RAM_35 = 256'hDCFF90043000039300D000FFF3FB38FE5F0035C9EC000243FFC3E60BF5FBC801;
defparam prom_inst_16.INIT_RAM_36 = 256'hFEE182359EFFC00A6000072601A001FFFFFFF0FCFE009AD716003743FBE1D3E0;
defparam prom_inst_16.INIT_RAM_37 = 256'h74006E8FF8E4C25F9DE782164C000E4C034003FFF1F1F8FE5C000AAA9C011DF7;
defparam prom_inst_16.INIT_RAM_38 = 256'hD80004C3FBFE77FB06646C7819FF802D40003C98028007FFE3FFF8EEA86038DC;
defparam prom_inst_16.INIT_RAM_39 = 256'h0BE2E70DCC000C731E9FEFFF1716977ADDEE40AA8000793005000FFF87F48B84;
defparam prom_inst_16.INIT_RAM_3A = 256'h14003FFE16F9CF0BBD000E7B0F1FFFF8201325FADDFC9F350000F2600A001FFF;
defparam prom_inst_16.INIT_RAM_3B = 256'h0001C98028007FFC24EF9E162240263DA9FFFFF0201721EE99A819AE0001E4C0;
defparam prom_inst_16.INIT_RAM_3C = 256'hC5728ED8000393005000FFF80DF7E7AFD080619F8CEFF80200037CFBC130277C;
defparam prom_inst_16.INIT_RAM_3D = 256'h4302FCF80121999000072600A001FFF06FBF8FF21200000FC50FF0000003FCBB;
defparam prom_inst_16.INIT_RAM_3E = 256'hE004003002CBE705B4821320000E4C014003FFE0CF8D1E4538001867700380E0;
defparam prom_inst_16.INIT_RAM_3F = 256'hA7800703EC00AA1068F778C3030E7260003C9006CFFFFFC198DA3C7CAC001C24;

pROM prom_inst_17 (
    .DO({prom_inst_17_dout_w[30:0],prom_inst_17_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_17.READ_MODE = 1'b0;
defparam prom_inst_17.BIT_WIDTH = 1;
defparam prom_inst_17.RESET_MODE = "SYNC";
defparam prom_inst_17.INIT_RAM_00 = 256'hFFEF70EDE0000F01EB2869C1647E6003811CFCE00079200D900FFFFFFF165255;
defparam prom_inst_17.INIT_RAM_01 = 256'h003FFFFFF66E764A78201FF16740060FDF92607311AD31C000F24019001FFFFF;
defparam prom_inst_17.INIT_RAM_02 = 256'h03C90024007FFFFFEF7FD0334E4003C1ADFF8E5709B54057221C62C001E48032;
defparam prom_inst_17.INIT_RAM_03 = 256'h3EF32A000792006800FFFFFFFC7CF4A8188001901B72D310D43E00171C789580;
defparam prom_inst_17.INIT_RAM_04 = 256'h35520615FDBE14000F2400D001FFFFFFEFF9C6FF910000103BF457C6D95D0713;
defparam prom_inst_17.INIT_RAM_05 = 256'h162604AE007B0607E63038001E4801A003FFFFFED9F2CF85E800001E7D1DCF93;
defparam prom_inst_17.INIT_RAM_06 = 256'hA64606059C5A354B7FB40600F24120003890036007FFFC0136704EA384000001;
defparam prom_inst_17.INIT_RAM_07 = 256'hE5DF0513FF04BE0057BBD3CB65AB8E0CE7C26000712006800FFFFF01F66F82EC;
defparam prom_inst_17.INIT_RAM_08 = 256'h3FFFF8036AFF1FCBEF02FFEF583FAB6E88800E0999C5C000E2400D001FFFFC03;
defparam prom_inst_17.INIT_RAM_09 = 256'hC90024007FFFE0027DBFF5CC04401FFF13E2667360C31E09229AC001E4801A00;
defparam prom_inst_17.INIT_RAM_0A = 256'hFA5900079200C800FFFF8004CE7FF505A8803FFD0DB6B1F5D2C00F0A7EB48003;
defparam prom_inst_17.INIT_RAM_0B = 256'h89133F17D9F0000F24019001FFFF000F967F8D0183E53F7FC42A6C1628839F12;
defparam prom_inst_17.INIT_RAM_0C = 256'h5CDE38265D55D81486E0001E48032003FFFE000DCE7EB680A2327FFD2847009F;
defparam prom_inst_17.INIT_RAM_0D = 256'hCBB9FFFE07253B2CCC27825F8B00087CD0028007FFFC004B58FFD0805420FDFA;
defparam prom_inst_17.INIT_RAM_0E = 256'hD8FF08097FBFF3EE2138FD3644A58E2EBE0000F9A005000FFFF800123C7F84C6;
defparam prom_inst_17.INIT_RAM_0F = 256'hFF80006219FF0C1E499FE7DE150FC8C2FB8F3C57F80001F3400A001FFFE00031;
defparam prom_inst_17.INIT_RAM_10 = 256'h006A007FFE00005AB3FF11295C3FF1FFA4D86D212777DDE9D00003E68014003F;
defparam prom_inst_17.INIT_RAM_11 = 256'h18000F9A00D600FFF0000033FBFF0690AE1FE1CF2BB1E7BE878F97324C0007CD;
defparam prom_inst_17.INIT_RAM_12 = 256'hF947EE1834001F3401AC01FFC0000065F3FF704B780F1F1FBE88217B06FFA7C6;
defparam prom_inst_17.INIT_RAM_13 = 256'hFC0FA1646880F67068003E68035803FF0000014DE7FF31CF50060E1F224D74C1;
defparam prom_inst_17.INIT_RAM_14 = 256'h80020816EE428CCA80FD0BF9E0003CD006B007FC000002C3C7FC86C4F0030C47;
defparam prom_inst_17.INIT_RAM_15 = 256'hBDFD888F400609AD47CE9C388FE5E363800079A00D600FFF87000EE73EFED70C;
defparam prom_inst_17.INIT_RAM_16 = 256'h001FFD2B3FFB9801E00E107A18C2283443B37DCF8000F3401AC01FFF0000FFDC;
defparam prom_inst_17.INIT_RAM_17 = 256'h6B007FE003FFFC977FF6344BC00C401778D83D324CE17ABF0001E68035803FFC;
defparam prom_inst_17.INIT_RAM_18 = 256'h00079A10D600FFFF7FFF898E7FFC6AF7001CE02E17447DFB959EF27E0003CD00;
defparam prom_inst_17.INIT_RAM_19 = 256'h689287FE000F3421AE01FFFFFFFF01CEFFF483CE00387143E7DDDBB8139AD3FF;
defparam prom_inst_17.INIT_RAM_1A = 256'h9E5534B20F18FFFC001E68635C03FFFFFFF0115CFFE9433C007078C70E618734;
defparam prom_inst_17.INIT_RAM_1B = 256'h03E5713653B511884F6DD038003CD3C6B007FFFFFF802399FFC03AF801FC3D3F;
defparam prom_inst_17.INIT_RAM_1C = 256'h3FCC64F00780393C02D6D1B4D5AC9F700079A78D600FF87BF00420BF9FDC36E0;
defparam prom_inst_17.INIT_RAM_1D = 256'h0004847F7F68E7800E38A7602B78E717DD383EE000F34F1AC01FF1FFC000413F;
defparam prom_inst_17.INIT_RAM_1E = 256'h00403FFC00DC967EEB9128003CC06D454FA7D164277A5DC001E69E35803FFFFF;
defparam prom_inst_17.INIT_RAM_1F = 256'h079E78D600007FF81FB905FF99B1F6007FDEDC99FBB625883AA41F8003CD3C6B;
defparam prom_inst_17.INIT_RAM_20 = 256'h5B5C3C000F3CF1BC0003FFFEFF7317DF3685B8F8CC61FC1102A4577068723F00;
defparam prom_inst_17.INIT_RAM_21 = 256'h062017608E2D78001E79E378000FFFFFFFC63FBE7D158FF9045A5B13BC4C6410;
defparam prom_inst_17.INIT_RAM_22 = 256'h5F7469485F90896190DC27B01CD1C670003FFFFFFF182F3C714913FA93905972;
defparam prom_inst_17.INIT_RAM_23 = 256'h61CA133BB9E6666AB2E09522286DE50079A78CE000FFFFFFFFE04F35F8C1DDC1;
defparam prom_inst_17.INIT_RAM_24 = 256'hFFD85ED683F3647605D79B4F4971946EFC388A00F34F1958007FFFFFFFC0EE6A;
defparam prom_inst_17.INIT_RAM_25 = 256'h00FFFFFFFFF3BDEE07F87AAC1053968C9150E0A0655C3D81E69E32FC001FFFFF;
defparam prom_inst_17.INIT_RAM_26 = 256'h9AF8C9F000FFFFFFFFE63FCC833FA29DFA875611FBE923731910BC83CD7C65FC;
defparam prom_inst_17.INIT_RAM_27 = 256'h5365360735F993C0381FFFFFFF697FD956253CB3E3C85E5CBF7517EF47A03003;
defparam prom_inst_17.INIT_RAM_28 = 256'h2034AF8372D190066BF30601981FFFFFFEC6FFEEBD614D4EC10BBA87A3C504C0;
defparam prom_inst_17.INIT_RAM_29 = 256'h76AC399D57E14022FCF98D8F57C61F04803FFFFFFD91FFDF7837DC9CE3C6886F;
defparam prom_inst_17.INIT_RAM_2A = 256'h6DA1307A3DDB04D6A7C3A06320CBE50EAF8C3E0F200BFFFFFBA4B5493688883F;
defparam prom_inst_17.INIT_RAM_2B = 256'hFE3D56A6D06170D4B7A615E48CC8E300B7105A1D5F1C3C1F3013FFFFF707EA52;
defparam prom_inst_17.INIT_RAM_2C = 256'hE807FFFFFC12AF0D9D14E02FC27F2C63698A46282804843ABE38783F9807FFFF;
defparam prom_inst_17.INIT_RAM_2D = 256'hF8F4F8FE6807FFFFD82DC71B883560507FFF3D695E12972B015640F57C72F84F;
defparam prom_inst_17.INIT_RAM_2E = 256'h6DED23D5F1E9FFFC1807FFFFF8CB06B7F2D3C0A0303E7D723868EE2D44BB01EA;
defparam prom_inst_17.INIT_RAM_2F = 256'h2620F1F9EED95FABE3D0FFF81407FFFFF19AA56EE317A060827CEE2132B5E563;
defparam prom_inst_17.INIT_RAM_30 = 256'hC0E582AC926E5C033F2F5427E7B7FDE01807FFFFD0B54AD647B1409184F8BBA9;
defparam prom_inst_17.INIT_RAM_31 = 256'h10641F17C1CB8B5CA708E66DD1EFC84FCF6FF1C03007FFFE622B85F7C83A0F99;
defparam prom_inst_17.INIT_RAM_32 = 256'hC4E357F860C82E3F83972DC71239497F933E309F1EC1E180780FFFFE44770BEC;
defparam prom_inst_17.INIT_RAM_33 = 256'h26DFFFFC8146AFF0E5840C3F0E0ED06C3494F00CBEB8613E3F80C000EA3FFFFE;
defparam prom_inst_17.INIT_RAM_34 = 256'hBE000000348FFFF9189C7F61EBDC1C3C1C1DF0206172F356E300C37C5F000000;
defparam prom_inst_17.INIT_RAM_35 = 256'hAFAF0CE17C020000410FFFF35358DA63DDBC1800783BC1B8FEC5A2CB916186F8;
defparam prom_inst_17.INIT_RAM_36 = 256'hD6A7ECD5B34239C2F80C7810E00FFFE6973DB2C7B9783001E062E82753825EE8;
defparam prom_inst_17.INIT_RAM_37 = 256'h83A6CC093E338A7F5A203705D818F020901FFFBD6E79648772F07003C0877979;
defparam prom_inst_17.INIT_RAM_38 = 256'hE785C0FF074C716935B5B85311DA6E0BB030062080FFFFF905BC641E75C2C87F;
defparam prom_inst_17.INIT_RAM_39 = 256'h86319C7EC40FC3FE0E826144DE193BB57FA0DC1660600C0141FFFFFAC718C23E;
defparam prom_inst_17.INIT_RAM_3A = 256'h07FFFFE63D030474C81F8FF83D00CFF47DE82EFD8BA7382CC1C0180183FFFFF4;
defparam prom_inst_17.INIT_RAM_3B = 256'h070000450FFFFFC8500738A5F03FBFF07B007187992230470856F05D83802022;
defparam prom_inst_17.INIT_RAM_3C = 256'hA40DC10E0E0000841FFFFF568D0E40D0746FFFE0F65C6C4831EE526CB774E0BF;
defparam prom_inst_17.INIT_RAM_3D = 256'h2DB1D7D16217831C1DFE700A1FFFFEB4025C51D7269BFFC1E5134C62F3003E5C;
defparam prom_inst_17.INIT_RAM_3E = 256'hD62ADB76FBBD14360C2602C10BFCE0143FFFFD3194BAE38E5937FF03CF713FAB;
defparam prom_inst_17.INIT_RAM_3F = 256'h8FFFF80FACD1E01BDAD31FE7384E05801FFFF8929FFFFFDCCCBCC7B71BFFFC07;

pROM prom_inst_18 (
    .DO({prom_inst_18_dout_w[30:0],prom_inst_18_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_18.READ_MODE = 1'b0;
defparam prom_inst_18.BIT_WIDTH = 1;
defparam prom_inst_18.RESET_MODE = "SYNC";
defparam prom_inst_18.INIT_RAM_00 = 256'h92ED8F021FDFF01751B4017588F08E02509C1A203FFFF1253FFFFFA8197F861D;
defparam prom_inst_18.INIT_RAM_01 = 256'hFFFFFFBC63591D6B3FFF800E837B3B8EC3B536C1A13834403FFFE2427FFFFF1E;
defparam prom_inst_18.INIT_RAM_02 = 256'hFFFF81C1FFFFFECCC4E21A5FFFFC001D05B274F436D0DAB9C27068807FFFC0A0;
defparam prom_inst_18.INIT_RAM_03 = 256'h09C0B001FFFF6382FFFFF88989D810DBFFF0003A4A787B7924A5DE7784E0D100;
defparam prom_inst_18.INIT_RAM_04 = 256'hA977FEB613816203FFFEC745FFFFF0C333722993FFC0006C95D0FF3EDA1472D3;
defparam prom_inst_18.INIT_RAM_05 = 256'h8EE7CA72132D30303F82C87FFFFD848BFFFFE3C2F6D42C87C38005995B2706AD;
defparam prom_inst_18.INIT_RAM_06 = 256'hF510369D1D4B18142DFA016D9F05D1FFFFFE0937FFFFE6178B885300E3400B4A;
defparam prom_inst_18.INIT_RAM_07 = 256'h1FC6AEE1E260FD7AB106C19DD2335638BE0FA7FFFFFC126FFFFFC0235F10199F;
defparam prom_inst_18.INIT_RAM_08 = 256'hFFFFC808B38E000FF3C1F2FD40B35E190B2EDDE1BC1DBFFFFFFB24DFFFFFC644;
defparam prom_inst_18.INIT_RAM_09 = 256'hFFFE117FFFFFF043E71CAB07C387ED7BA1A567AE33FA100BFC3B7FFFFFFF08BF;
defparam prom_inst_18.INIT_RAM_0A = 256'hF1BDFEFFFFFEE2FFFFFFEA87CEBE9900821F9EE773E51F04A757BEA4F856FFFF;
defparam prom_inst_18.INIT_RAM_0B = 256'hAC696C17E37BFC07FFFDC5FFFFFFF46DBC2E0838E07F2DCFF6B1F6C851C022A5;
defparam prom_inst_18.INIT_RAM_0C = 256'hCED4FDA7320F8827E6F7F803FFFB8BFFFFFFF8FBF8EE80F280FE519FAF6061A9;
defparam prom_inst_18.INIT_RAM_0D = 256'h07CC8FFF9E40E922AE13504FCDAFF81FFFFD81FFFFF4F51FF24EC78003F1D7FF;
defparam prom_inst_18.INIT_RAM_0E = 256'hC5DFFE001F313FFF3D80A9861864009F9A1FFFFFFFFB03FFFFE9EA3FE06F0000;
defparam prom_inst_18.INIT_RAM_0F = 256'hFFA788FFE8FE47003EC6FFFE78D05E7D74F2C13F247FFFFFFFF607FFFFD3C47F;
defparam prom_inst_18.INIT_RAM_10 = 256'hFFBC0FFFFF4C11FFDFF88780396D7FFCBFB911FCE945027E48FFC7FFFFDC07FF;
defparam prom_inst_18.INIT_RAM_11 = 256'h23FEFCFFFF781FFFFE88B5FFF7C00781CD9FFEF97E513E94926D04FC91FF7FFF;
defparam prom_inst_18.INIT_RAM_12 = 256'h87EC13625FFE01FFFFF03FFFFD016AEFE3801F07252FF9F307F93B7728C209B9;
defparam prom_inst_18.INIT_RAM_13 = 256'hFE8EEF743EC22666971CC7FFFFF07FFFF802D5DE73C03F0EB2DBF3E47F831326;
defparam prom_inst_18.INIT_RAM_14 = 256'hC3FE7F007335B51B6EC30C0D6037D1FFFEC07FFF0D8BD69FF1F8C7C679FF3F81;
defparam prom_inst_18.INIT_RAM_15 = 256'h5F0783E307FCFE0249A527068CE0B80DE0E261FFF990FFC0CB17A7FFD8F1CECF;
defparam prom_inst_18.INIT_RAM_16 = 256'hE85E9FFCB81FF00D9FFFFC6CD8DD9D2CD423A02847F02B7FF721F01FD62F5E6E;
defparam prom_inst_18.INIT_RAM_17 = 256'hFC007FE7E0BCB56F13FF83B9FFFFFA8813BCC5DDB18E40509FBDA9BFE600C1FD;
defparam prom_inst_18.INIT_RAM_18 = 256'hECF85BF8F7FF00FF41799BBC67FF001AFFFFFD3924DCBF5B4FCC80B13C597DFF;
defparam prom_inst_18.INIT_RAM_19 = 256'h87CE03B72EDC7BE1F3800EE0A2F22646EE0007F5F7FFFAD1D9C372A9E48B01B3;
defparam prom_inst_18.INIT_RAM_1A = 256'hD180908842480FA1478CB780A0003C1145E41747D0003DEBEFFFF6C81F3D48CA;
defparam prom_inst_18.INIT_RAM_1B = 256'h3FFF97C3747144DE06C01F5D0F869B728DC7C00A457E780F8C081FD79FEFC557;
defparam prom_inst_18.INIT_RAM_1C = 256'h38003C583FFF2C5A9F9D1AE000D03EA41F8836ED3B1F00748649C03F1C003F2E;
defparam prom_inst_18.INIT_RAM_1D = 256'h124C81F878003CB47BFE2F90070943B0D5601D943FCBE9FE507C03EB228D00FE;
defparam prom_inst_18.INIT_RAM_1E = 256'h3F00FF961C7707F0F0007DF0F3FC426FE5DD713DBCC439DC79DCA3E313C01FC7;
defparam prom_inst_18.INIT_RAM_1F = 256'hE1FA2FD876007FBC74D81FC1F000F881E7FD93130FDE523938C8F87B71DEE7E0;
defparam prom_inst_18.INIT_RAM_20 = 256'h2373FDDCE9FADFC8E0003F3B57E27F03E001F1D7CFFAF1C7DEC2CD33D9B9F5FA;
defparam prom_inst_18.INIT_RAM_21 = 256'h5C12AA6766E609E1D87ABFB1C0003E751F30FC07C001E7AF9FE2EA5BB248D670;
defparam prom_inst_18.INIT_RAM_22 = 256'hC58F17681858F127FDCC1120CCF83B01E001FC574703E01FC005C5FF632FB1AD;
defparam prom_inst_18.INIT_RAM_23 = 256'h0003105FBF13102FA86542623B9827A1D9F17EB3C003F8ABBE07C03F80098BAE;
defparam prom_inst_18.INIT_RAM_24 = 256'hF83F01FC000601BFEF0F6D136D42AE81BF300E4390FC3C978007F2DC5C0F80FF;
defparam prom_inst_18.INIT_RAM_25 = 256'h001FCA3DF07C07F80004227FFE2C95AAA503BEB27E600603C066FECD000FE718;
defparam prom_inst_18.INIT_RAM_26 = 256'h11EBF16D003FD17FE0F80FF0004A69FFF06ED5C6AC65DDA1FCC00C0380F9FC4F;
defparam prom_inst_18.INIT_RAM_27 = 256'hF340CC063353E31A007FA2BFC1F03FE00094F7FFA32D388F78123FB3F9806003;
defparam prom_inst_18.INIT_RAM_28 = 256'hA5281D2EE5F18C266FF3EFB400FC561B83E07F80012967FF44885F39F01297FB;
defparam prom_inst_18.INIT_RAM_29 = 256'h3C41C4A1CD78048DCBE39E0ECC07CEF8000173FE0780FC00045FFA7AAE753A23;
defparam prom_inst_18.INIT_RAM_2A = 256'h1153E7FBF0B225528EFF14DB97C53C0FD48FDC70001E7BFC0F03F00008BFF4FF;
defparam prom_inst_18.INIT_RAM_2B = 256'h3C0FC0000322AFD34BF512169CCF29372E8A7C0D8BEFB8C0007867781E07E000;
defparam prom_inst_18.INIT_RAM_2C = 256'h03F3FF40F03F800006E56FCC6C5B6D33578FE06E4014F819074F39C001F1AEB0;
defparam prom_inst_18.INIT_RAM_2D = 256'h073CC0000FE69E01E0FF000005EB5F5D7CBA9227CDC755DC8014F838065E7380;
defparam prom_inst_18.INIT_RAM_2E = 256'h0152F028467AA0001FE1FA07C1FE0000414EB6F44552923FF4C6EBB80029F838;
defparam prom_inst_18.INIT_RAM_2F = 256'hCDC43ECAD304F05184F6A0003C4FF40F07FC0000811CEDDDECE9753E4C83F370;
defparam prom_inst_18.INIT_RAM_30 = 256'hD8C00FCDA4B34C918601FC93B3E41077057FF41C0FF800001FDD67FBED58E78A;
defparam prom_inst_18.INIT_RAM_31 = 256'h75BAC7D4DE1CEF9BCF0499220C0FF0B701D930CC757FE8701FF000003DDAC7F3;
defparam prom_inst_18.INIT_RAM_32 = 256'hFF0000004B758F3F093E0D77B64930451C3C68B7B1B3F003137F90E07FC00000;
defparam prom_inst_18.INIT_RAM_33 = 256'h21FE0F83FE0000007DE58E434BF0827F0DDEE096A848D137BB8BF0F3927F01C0;
defparam prom_inst_18.INIT_RAM_34 = 256'h777F4E07FFF81E07F80000003FE901D936508CEF1DEDC12910D1E1258783CC7C;
defparam prom_inst_18.INIT_RAM_35 = 256'h03A1F1B2CF46861FFFF07C1FF0000100A7E8068FB2D7FF4D1FFB82C20191F078;
defparam prom_inst_18.INIT_RAM_36 = 256'hBE9FCB9E7F63F7146CCD9C72BFE0F83FE000020027D20C59D47FFEC91B930584;
defparam prom_inst_18.INIT_RAM_37 = 256'h7F634FEAECBF94B17E47E2227B983380BF81E07F0004000177D400281DDB3BD7;
defparam prom_inst_18.INIT_RAM_38 = 256'h478C00EABF679BC7993F29E79C87E20F7E004E02FF03C0FE000800010E45D13B;
defparam prom_inst_18.INIT_RAM_39 = 256'h00200022116C09D87722A3F5357E43DBD3A4621BA0E13C09FE0783FC00100000;
defparam prom_inst_18.INIT_RAM_3A = 256'hF0781FE001C0004E1FCC909E7344476AB8FC9FA3074C4410E83CF017783E07F8;
defparam prom_inst_18.INIT_RAM_3B = 256'hEFFF00BDC0F07F800780001EC8C822BF745A0A7C21F9BB720648445C21838076;
defparam prom_inst_18.INIT_RAM_3C = 256'h0818C75163FE033F81E1FF001F00003FA5D0038E2C66F4FA03F370472C98461D;
defparam prom_inst_18.INIT_RAM_3D = 256'hCFDC46565094B445FB000ECE0383FC007E00000628E50246F3CBEAF467E7E202;
defparam prom_inst_18.INIT_RAM_3E = 256'h4996FFE80FB81D26D3884473780019D83F0FF807F80000393B075F8E69DBB7F7;
defparam prom_inst_18.INIT_RAM_3F = 256'hE6C67CEA146D7FD85F70F67DA720CCFE630833B07E1FF00FF000003719C1BE9D;

pROM prom_inst_19 (
    .DO({prom_inst_19_dout_w[30:0],prom_inst_19_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_19.READ_MODE = 1'b0;
defparam prom_inst_19.BIT_WIDTH = 1;
defparam prom_inst_19.RESET_MODE = "SYNC";
defparam prom_inst_19.INIT_RAM_00 = 256'hC000003FE2A4349518077FB5FEEFA1FF2F304C9E6FD0C7E0FC3FE01FE000003F;
defparam prom_inst_19.INIT_RAM_01 = 256'hE07FFFFF8000007FE2D93F7321A8FF7CFDC447FF2F008F60FFE18F01F83FFFFF;
defparam prom_inst_19.INIT_RAM_02 = 256'hFF062C0F00FFFFFF0000007F848249BD0ADCFE39FBB43F7F4F61E661FFC33607;
defparam prom_inst_19.INIT_RAM_03 = 256'h5E4EF9FFFE1CD01E01FFFFFE000001FF848C4EB99D71FD73F7487F3F4F43C4E1;
defparam prom_inst_19.INIT_RAM_04 = 256'hDD83777E9EDDFA1FF8F9203C03FFFFFC000003FF8C8D5CB5B833F9AFEE82EF3F;
defparam prom_inst_19.INIT_RAM_05 = 256'h0000000000000166B6FE3A1C31EFC07807FFFFF800003BFF1E34139440C4C8DF;
defparam prom_inst_19.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_19.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_20 (
    .DO({prom_inst_20_dout_w[30:0],prom_inst_20_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_20.READ_MODE = 1'b0;
defparam prom_inst_20.BIT_WIDTH = 1;
defparam prom_inst_20.RESET_MODE = "SYNC";
defparam prom_inst_20.INIT_RAM_00 = 256'hF010F4F7FFFFFFE010000000C3FFE0000000000000000003FFFFFCC7F8087AF5;
defparam prom_inst_20.INIT_RAM_01 = 256'hFFFFF31FE0206DFFFFFFFFC02000000187FF80000000000000000007FFFFF98F;
defparam prom_inst_20.INIT_RAM_02 = 256'h0000003FFFFFE63FC00001FFFFFFFFC0400000021FFF0000000000000000001F;
defparam prom_inst_20.INIT_RAM_03 = 256'h000000000000007FFFFF8C7FC0006D1FFFFFFE81800000003FFE000000000000;
defparam prom_inst_20.INIT_RAM_04 = 256'hFFF0008000000000000000FFFFFF08FFC000EC1FFFFFFA02000000007FF80000;
defparam prom_inst_20.INIT_RAM_05 = 256'h0001F1C3FFE0018000000000000001FFFFFE19FF8001E81FFFFFF80800000021;
defparam prom_inst_20.INIT_RAM_06 = 256'hFFFFC0400003FF8FFFC0030000000000000003FFFFFC31FF0003EC3FFFFFD020;
defparam prom_inst_20.INIT_RAM_07 = 256'h000FF237FFFE01000007F81FFFE7E60000000000000007FFFFF8C7FF0007FC7F;
defparam prom_inst_20.INIT_RAM_08 = 256'hFFE31FFC001FEC1FFFFA0200000FF03FFFCFCC000000000000000FFFFFF18FFE;
defparam prom_inst_20.INIT_RAM_09 = 256'h0000FFFFFFC63FFE003FF82FFFF00800001FE07FFF9F98001800000000001FFF;
defparam prom_inst_20.INIT_RAM_0A = 256'h7FFF80000003FFFFFF843FFF607FF01FFFD03000003FC1FFFF3F30003C3C0000;
defparam prom_inst_20.INIT_RAM_0B = 256'hFCFCC003FFFF0000010FFFFFFF083FFEE0FFF03FBFC04000001F83FFFE7E6000;
defparam prom_inst_20.INIT_RAM_0C = 256'h00020FFFF9F9800FFFFE0000063FFFFFFE107FFDE1FFF17F7E018000000707FF;
defparam prom_inst_20.INIT_RAM_0D = 256'hF0C0080000001FFFF3F3003FFFFC00001CFFFFFFFC207FFBC3FFF67FFA420000;
defparam prom_inst_20.INIT_RAM_0E = 256'hCFFFF87FC310000006003FFFC70383FFFFF80039FFFFFFFFF86007FFE7FFF4FF;
defparam prom_inst_20.INIT_RAM_0F = 256'hE19FFFFFDFFFF4FFD840000008007FFFCE0F03EFFFC00071FFFFFFFFF0CFFFFF;
defparam prom_inst_20.INIT_RAM_10 = 256'hFFFFFFFFC33FC0FFFFEFF5FE308000000000FFFFFC07FFFF9FFC00E1FFFFFFFF;
defparam prom_inst_20.INIT_RAM_11 = 256'h80000381FFFFFFFF867F80FFFFFFF5FE220000000001FFFFF8070FF83FFC01C1;
defparam prom_inst_20.INIT_RAM_12 = 256'hE0FFCFFF00000700FFFFFFFF0CFF00FFFFFFF7F00C0000000003FFFFF07FFCFF;
defparam prom_inst_20.INIT_RAM_13 = 256'h000FFFFFC0FDCFFFC0020E01FFFFFFFE19FE01FFFFFFF5D5100000000007FFFF;
defparam prom_inst_20.INIT_RAM_14 = 256'h80000000001FFFFF83EC7FFF00041C03FFFFFFFC33FC03FFFFFFF7DE40000000;
defparam prom_inst_20.INIT_RAM_15 = 256'hFFFFE2D200000000003FFFFC3F7FFFFC0007FEB7FFFFFFE047F803E7FFFFFE68;
defparam prom_inst_20.INIT_RAM_16 = 256'h9FE1C7FFFFFFF3A400000000007FFFF7FD0FFFF00010356FFFFFFFC08FF0C7EF;
defparam prom_inst_20.INIT_RAM_17 = 256'hFFFFFE033FE38FFFFFFFCD100000000000FFFFFFE81FFFE00030059FFFFFFF01;
defparam prom_inst_20.INIT_RAM_18 = 256'h019FFFFFFFFFB8067FC58FFFFFFFA8400000000001FFFFFF01FFFFC000F8033F;
defparam prom_inst_20.INIT_RAM_19 = 256'hC7FFFE0003FFF3FFFFFFF80CFF890FFFFFFFC8800000000003FFFFFF01FFFF80;
defparam prom_inst_20.INIT_RAM_1A = 256'h0FFFFFE21FFFF80007FFAFFFFFFFF019FF111EFFFFFF0A000000000007FFFFD4;
defparam prom_inst_20.INIT_RAM_1B = 256'h000000001FFFFD8807FFF0000DFBDBFFFFFFF033FE233DFFFFFF840000000000;
defparam prom_inst_20.INIT_RAM_1C = 256'hFFFFE000000004003FFECE0006FFE00007FFDFFFFFFFC063F8423DBFFFFFD800;
defparam prom_inst_20.INIT_RAM_1D = 256'hE106673FFFFF80000000F8007FFF61E83FFF80000FFF3FFFFFFF80C7F0867F9F;
defparam prom_inst_20.INIT_RAM_1E = 256'hFFFE031FC204E73FFFFF98000001F000FFF4B05E0FFF0001FFFF3FFFFFFF018F;
defparam prom_inst_20.INIT_RAM_1F = 256'hFFFEFFFFFFFC063FC40CC67FFFFED0000006C001FFD4001F1FFE0007FFFE7FFF;
defparam prom_inst_20.INIT_RAM_20 = 256'hF7F8000FFFFFFFFFFFF80C7F8808967FFFFF500000188003FF6A000FFFFC000F;
defparam prom_inst_20.INIT_RAM_21 = 256'hF0100001FFF0001FFFFFFFFFFFF018FF101814FFFFFF200000210007FC1B0007;
defparam prom_inst_20.INIT_RAM_22 = 256'h0374001DE04000017FE0001FFFFFFFFFFFE031FE2010107FFFFF200001DA000F;
defparam prom_inst_20.INIT_RAM_23 = 256'hFFFE000006E8003301600001BF800077FFFEEFFFFFC067F8461090FFFDFEC000;
defparam prom_inst_20.INIT_RAM_24 = 256'h003031FFFFFF000019D0006002000000CE0000EFFFFDFFFFFF80CFF0843010FF;
defparam prom_inst_20.INIT_RAM_25 = 256'hFE031FC2003016FFFFFD000077A000C148000000CC0000FFFFFCFFFFFF019FE1;
defparam prom_inst_20.INIT_RAM_26 = 256'hFFF9FFFFFC063F84006017FFFFFC0000DF4001804000000C4600007FFFFDFFFF;
defparam prom_inst_20.INIT_RAM_27 = 256'h2800003FFFF1FFFFF80C7F0800E037FFFFFE00033E80031080000000400000BF;
defparam prom_inst_20.INIT_RAM_28 = 256'h000006E0F400007FFFF3FFFFF018FE1001E02FFFFFF00004FD000C7400000000;
defparam prom_inst_20.INIT_RAM_29 = 256'hEC00306800000F39F400007FFFAFFFFFE031FC2013E02FFFFFF8001BF20018A0;
defparam prom_inst_20.INIT_RAM_2A = 256'hFBFC8197E8026440000003DF7FC000FFFF8FBFFFC067F8C007E02FFFFFFC006F;
defparam prom_inst_20.INIT_RAM_2B = 256'h0F005FFFFFF3C0FFB000D700000003EFFF0001FFFF2FFFFF80CFF1800F80BFFF;
defparam prom_inst_20.INIT_RAM_2C = 256'h033FC6001E005FFFFFF0023F60012400000003EFFBE300FFFEDFFFFF019FE300;
defparam prom_inst_20.INIT_RAM_2D = 256'hFF7FFFFC067F8C0003C05FFFFFFE213EC0077800000023DFFBE401FFFF9FFFFE;
defparam prom_inst_20.INIT_RAM_2E = 256'hFBC1E1FFFC5FFFF80CFF180007E07FFFFF9FB0BF800F800000000FFFFBC083FF;
defparam prom_inst_20.INIT_RAM_2F = 256'h001FCFFFFDE1F9FFF83FFFF019FE30000FC0BFFFFF60614D0009C00000009FFF;
defparam prom_inst_20.INIT_RAM_30 = 256'h00440000003FEFFEFFF8FFFFD0FFFFE033FC60001E00BFFFFF801BDA00118000;
defparam prom_inst_20.INIT_RAM_31 = 256'hFB801C6408E80000107FFFFFFDC4EBFFABFFFFC067F8EFE03C027FFDFD001A94;
defparam prom_inst_20.INIT_RAM_32 = 256'h0381FFFFF7000CC82080030041FFFFF779C1FFFF53FFFF80CFF1DFF001C47FFF;
defparam prom_inst_20.INIT_RAM_33 = 256'h3FC7FFC00700FFFFE8000D38000013C00FFFFFF329D3FFFF87FFFF019FE3FFE0;
defparam prom_inst_20.INIT_RAM_34 = 256'h47FFFE067F8FFF800E03FFFFB0000622480023C07FFEFFF80DFFFFFF8FFFFF03;
defparam prom_inst_20.INIT_RAM_35 = 256'h00FFFFFC8FFFFC08FF1FFF000C01FFFFA0000710000003C3FFFFFFF009FBFFFF;
defparam prom_inst_20.INIT_RAM_36 = 256'hFFFFFFC800FFFFF95FFFF811FE3FFE000005FFFF80000318460037C3FFFFEF99;
defparam prom_inst_20.INIT_RAM_37 = 256'h7C007EFFFFFBFDE001FFFFF23FFFF023FC7FFC000E05FFFE2000028C9C011DF7;
defparam prom_inst_20.INIT_RAM_38 = 256'h000000C3FFFE77FBFFFBF38001FFFFE43FFFC047FCFFF8001C0BFFFE400000CA;
defparam prom_inst_20.INIT_RAM_39 = 256'hF40BFFF20C000073FEFFEFFFFFF9F88201EFFF987FFF808FF9FFF0007800FFF9;
defparam prom_inst_20.INIT_RAM_3A = 256'hE7FFC001E817FFF43C00007BFFFFFFFFFFFCF80201FFFF10FFFF011FF3FFE000;
defparam prom_inst_20.INIT_RAM_3B = 256'hFFFE047FCFFF8003D81FFFE03800203DDFFFFFFFFFF8D81601EFF861FFFE023F;
defparam prom_inst_20.INIT_RAM_3C = 256'h01FD81C7FFFC08FF9FFF0007F027FFC3E800601FFFFFFFFDFFFC800301FFE0E3;
defparam prom_inst_20.INIT_RAM_3D = 256'hBCFC000201FF87AFFFF811FF3FFE000F902FFFA0E800000FFBFFFFFFFFFC0003;
defparam prom_inst_20.INIT_RAM_3E = 256'hFFFFFFCFFF340007317E0F5FFFF023FE7FFC001F302FFFA0C80018074FFFFF1F;
defparam prom_inst_20.INIT_RAM_3F = 256'hD0000703F3FF75E7970D000301FC0E1FFFC04FF8F000003E615FFFD9D8001C07;

pROM prom_inst_21 (
    .DO({prom_inst_21_dout_w[30:0],prom_inst_21_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_21.READ_MODE = 1'b0;
defparam prom_inst_21.BIT_WIDTH = 1;
defparam prom_inst_21.RESET_MODE = "SYNC";
defparam prom_inst_21.INIT_RAM_00 = 256'h00BFFFA200000F01E4D79E368380000381F81C1FFF809FF1EFF00000005FDF0C;
defparam prom_inst_21.INIT_RAM_01 = 256'hFFC0000000FFFD9980001FF1E83FF9F1C06C00031160F03FFF013FE1FFE00000;
defparam prom_inst_21.INIT_RAM_02 = 256'hFC04FFC7FF800000017FFEEE800003C1E80071AC2FC900072383E03FFE027FC3;
defparam prom_inst_21.INIT_RAM_03 = 256'h3E0F01FFF809FF8FFF000000017FE972C00001907CCD4C7E6C6000071F07807F;
defparam prom_inst_21.INIT_RAM_04 = 256'h0C400607FC0E03FFF013FF1FFE00000002FFFFA1400000105CAB1BDC38C10703;
defparam prom_inst_21.INIT_RAM_05 = 256'h2DFE6589FC630605FC1007FFE027FE3FFC00000103FFF4BAA000001E4CB9378B;
defparam prom_inst_21.INIT_RAM_06 = 256'h1402060424E824D27DC00607F3209FFFC04FFC7FF80003FE07FEFC9850000001;
defparam prom_inst_21.INIT_RAM_07 = 256'h0FFFF95C0204BE00657B3D88EDA38E0FE7401FFF809FF8FFF00000FE03FFFCB3;
defparam prom_inst_21.INIT_RAM_08 = 256'hC00007FC06FFE5CC1703FFEF7EDDD7EE78C00E0F84823FFF013FF1FFE00003FC;
defparam prom_inst_21.INIT_RAM_09 = 256'h04FFC7FF80001FFC1DFFFDF7D7001FFF3E3993F050431E0F00893FFE027FE3FF;
defparam prom_inst_21.INIT_RAM_0A = 256'h4A26FFF809FF0FFF00007FF80EFFFDF9EF803FFF0A686FFC49C00F0E16837FFC;
defparam prom_inst_21.INIT_RAM_0B = 256'h04733F1E388FFFF013FE1FFE0000FFF03FFFF1FE5CC53F7FDB70FAF622039F1E;
defparam prom_inst_21.INIT_RAM_0C = 256'h4FA2FAE616C5DC1FE11FFFE027FC3FFC0001FFF05FFFD8FF2DA27FFF382853FE;
defparam prom_inst_21.INIT_RAM_0D = 256'hD5D9FFFE14CBB9FC0087865340FFF7804FFCFFF80003FFB03BFFECFF36E0FFFE;
defparam prom_inst_21.INIT_RAM_0E = 256'h7FFFF67340FFFFFE34E6F0EE03E78E3781FFFF009FF9FFF00007FFE0BFFFFEF9;
defparam prom_inst_21.INIT_RAM_0F = 256'h007FFF837FFFF46EB29FFFFE1BA3E37E278F3C5F27FFFE013FF3FFE0001FFFC1;
defparam prom_inst_21.INIT_RAM_10 = 256'hFF8DFF8001FFFF9AFFFFFF42E63FFFFFBF886AFC8177DDB84FFFFC027FE7FFC0;
defparam prom_inst_21.INIT_RAM_11 = 256'hFFFFF009FF19FF000FFFFFB1FFFFFC83161FFFFF7911F63D058F9F303FFFF804;
defparam prom_inst_21.INIT_RAM_12 = 256'hE6C7FE85FFFFE013FE33FE003FFFFF65FFFFEC5D280FFFFFD83FF37802FFBF42;
defparam prom_inst_21.INIT_RAM_13 = 256'hCB7FC507C983F40BFFFFC027FC67FC00FFFFFE49FFFFF2C6F007FFFFC9FFCAC1;
defparam prom_inst_21.INIT_RAM_14 = 256'h8003FFF7923E3A4F8CDF3D07FFFFC04FF8CFF803FFFFFCCBFFFFE0ED7003FFA7;
defparam prom_inst_21.INIT_RAM_15 = 256'hFDFFD0E50007FE6F7639F43F9BE7FC3FFFFF809FF19FF00078FFF0C7FEFFF83A;
defparam prom_inst_21.INIT_RAM_16 = 256'hFFE0012FFFFFA9D4000FFFFE74BC887F3073FC3FFFFF013FE33FE000FFFF018F;
defparam prom_inst_21.INIT_RAM_17 = 256'h8CFF801FFC00001FFFFE47A8000FBFDCB4B79DF5CC22F97F3FFE027FC67FC003;
defparam prom_inst_21.INIT_RAM_18 = 256'hFFF809FF19FF00008000705FFFFC8D50001F1FB9F5B7BFFDFB9FF3FE7FFC04FF;
defparam prom_inst_21.INIT_RAM_19 = 256'hC9938FFFFFF013FE31FE00000000F0BFFFF91E80003F8F77F5027FBFD09BCFFF;
defparam prom_inst_21.INIT_RAM_1A = 256'hECA59E67DD1B7FFFFFE027FC63FC0000000FE0FFFFF37980007F86EF7CB8CF33;
defparam prom_inst_21.INIT_RAM_1B = 256'h03FE8FB7A857363DED4FDFFFFFC04FF8CFF80000007FC1FFFFF6F70001FFC36F;
defparam prom_inst_21.INIT_RAM_1C = 256'h3FB7DC0007FFC7BFFF4DBC3D8BAD3FFFFF809FF19FF000000FFBC1FF9FC9EA00;
defparam prom_inst_21.INIT_RAM_1D = 256'hFFFB05FF7FCFB0000FFF43EFE2DF3E1F7935BFFFFF013FE33FE000003FFF83FF;
defparam prom_inst_21.INIT_RAM_1E = 256'hFF800003FF2303FEEB9F40003FFE775BC09CFD7DD7725FFFFE027FC67FC00000;
defparam prom_inst_21.INIT_RAM_1F = 256'hF809FF19FF000007E0460FFF99BF50007FED26A5EAA0FFFF5DF95FFFFC04FF8C;
defparam prom_inst_21.INIT_RAM_20 = 256'h057C3FFFF013FE23FE000001008C17FF33FC68F8FF438E29F1A3F7DBB3BDBFFF;
defparam prom_inst_21.INIT_RAM_21 = 256'h847F7A496020BFFFE027FC47FC00000000382FFE67F31BF9F849292B137BC5DA;
defparam prom_inst_21.INIT_RAM_22 = 256'h9FDE972BFB7F763137733C4FE04FF88FF800000000E40FFCCDC5EBFB64715D43;
defparam prom_inst_21.INIT_RAM_23 = 256'hA7CB8F3C38FFE163E5FA6CEC14421AFF809FF11FF000000000185FF5D3C1FBC6;
defparam prom_inst_21.INIT_RAM_24 = 256'h0020FFD54FFFE838025FF94E07AAF5DB060025FF013FE227E00000000030BFEA;
defparam prom_inst_21.INIT_RAM_25 = 256'h800000000001FFE99FEC74301EDFF08FEF2FEBD65C40227E027FC403C0000000;
defparam prom_inst_21.INIT_RAM_26 = 256'h09FF100F000000000002FFC3BFE2F861C80E701B4EFFF6B95161837C04FF8803;
defparam prom_inst_21.INIT_RAM_27 = 256'h1FAE8BF813FE203E380000000083FF877FB120C3A0C2E25E9EFEFD7B38CF8FFC;
defparam prom_inst_21.INIT_RAM_28 = 256'hBFE7F1433C3DDFF827FC41FE180000000107FF1AFF50798FF305DC983FF5F8A1;
defparam prom_inst_21.INIT_RAM_29 = 256'h37343D942FFF9906D58DE7F0CFF880FF000000000203FE35FEE8711E81AB8C4B;
defparam prom_inst_21.INIT_RAM_2A = 256'hEC808479C1F800BDDFFF223CDB9457F19FF101FFC0000000040FFC49F771723F;
defparam prom_inst_21.INIT_RAM_2B = 256'h002DF0A7C0E318D3378018BE7FFF96BDBF12EFE33FE603FFC00000000817F853;
defparam prom_inst_21.INIT_RAM_2C = 256'hF0000000003BE14FA30230200000207A1FFC5E153C109FC67FCC07FFE0000000;
defparam prom_inst_21.INIT_RAM_2D = 256'hFF2407FE70000000207FCB9F780C404F8000347DBFF0CE6D6C437F0CFF9A07CF;
defparam prom_inst_21.INIT_RAM_2E = 256'hBD9FFC33FE4801FC1000000000FF9FBEF230809FCFC07674FFD57DF2CD99FE19;
defparam prom_inst_21.INIT_RAM_2F = 256'hFF0517742C29E067FC9003F818000000017FBF7DE0F1201FFF80F639FF84DDDB;
defparam prom_inst_21.INIT_RAM_30 = 256'hFF05EC9BFE939FAE9D50689FF93005E01000000021FF7EF241EA407FFF00EAE5;
defparam prom_inst_21.INIT_RAM_31 = 256'h0F0800FFFE0BD8D3FD7D7FEC53AFE13FF26001C03800000182FF7DFFC784007F;
defparam prom_inst_21.INIT_RAM_32 = 256'h03F8B7D81E1001FFFC17B5E5FED5FF1E30DFC27FE4C001807000000185FEFBFC;
defparam prom_inst_21.INIT_RAM_33 = 256'h360000030F796FB01C2403FFF00F6063D5CFFE2D313F84FFCB800000F2000001;
defparam prom_inst_21.INIT_RAM_34 = 256'h2E000000240000061EF2DF60189C03FFE01EE0EFBFF7FF97957F08FF97000000;
defparam prom_inst_21.INIT_RAM_35 = 256'h1E3423FE5C0000006000000C0FC59EE0313C07FF803DF1C7AFCFE3EAB07F11FF;
defparam prom_inst_21.INIT_RAM_36 = 256'hAA79E8F6DF1867FCB8000010C00000183E073FC062780FFE007A91BB639FDAAF;
defparam prom_inst_21.INIT_RAM_37 = 256'h03C3317796EFC0484F888FF978000020D00000407C0E7F80C4F00FFC00F581A0;
defparam prom_inst_21.INIT_RAM_38 = 256'h37843F000787915DB07F06C0D9E11FF2F0000020C000000038747A0119C23780;
defparam prom_inst_21.INIT_RAM_39 = 256'hF9D1F401640C3C000F1793B922FEA5822FC23FE5E00000018000000078E8F600;
defparam prom_inst_21.INIT_RAM_3A = 256'h00000002F2E3EC02881870003E2F7E5CA16E89C61F82FFCBC000000100000001;
defparam prom_inst_21.INIT_RAM_3B = 256'h0000004600000001CDC7E801703040007C5F2EF9626B344C2F6DFF9780000023;
defparam prom_inst_21.INIT_RAM_3C = 256'h7823FE2E0000008600000083978FD0127A600000F8FB2FB57EF9B2D87893FF2F;
defparam prom_inst_21.INIT_RAM_3D = 256'hFB52C6AADC4FFC5C0000000C0000010E2F5FF033C2840001F97C1E9CCE67E0B1;
defparam prom_inst_21.INIT_RAM_3E = 256'hEDEDDC9B0E0B0785709FFC800000001800000214CEBFA067D9080003F2BEB3E2;
defparam prom_inst_21.INIT_RAM_3F = 256'h0000000FDBDEFAD8754E1C9FC13FF9000000009A00000000FC3FC07B18000007;

pROM prom_inst_22 (
    .DO({prom_inst_22_dout_w[30:0],prom_inst_22_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_22.READ_MODE = 1'b0;
defparam prom_inst_22.BIT_WIDTH = 1;
defparam prom_inst_22.RESET_MODE = "SYNC";
defparam prom_inst_22.INIT_RAM_00 = 256'h50FF810F00200017B7B65E7D0CDE3473A27FE3200000013400000011F87F0198;
defparam prom_inst_22.INIT_RAM_01 = 256'h000000C1E17E037A0000000F6F7D0A322B687E5244FFC6400000026000000040;
defparam prom_inst_22.INIT_RAM_02 = 256'h0000018000000097C0FE06740000001EDDFE8F38F640DA9209FF8C80000000C0;
defparam prom_inst_22.INIT_RAM_03 = 256'h27FF2000000003000000002F81FE08CC0000003DFBFF181E2485A43413FF1900;
defparam prom_inst_22.INIT_RAM_04 = 256'h9502F4D04FFE4200000006400000019F03FA199C00000073F76D89F6D1047C74;
defparam prom_inst_22.INIT_RAM_05 = 256'h8FB8302350CDACD08FFC8878000006800000037A87FC1CF8000005E7CF9AD462;
defparam prom_inst_22.INIT_RAM_06 = 256'hFB0037271F73F1CDE3BA088DBFF911F000000D00000007F60FF8C00003000B97;
defparam prom_inst_22.INIT_RAM_07 = 256'h1FE2FF1E1E00FE0EBDFF03916ED1D4A27FF227E000001A00000003E85FF9E9FF;
defparam prom_inst_22.INIT_RAM_08 = 256'h00000320BFF01C0FF001FC1D7BFDA056F4EFDD2C7FE63FC000003400000001D0;
defparam prom_inst_22.INIT_RAM_09 = 256'h0000500000000641FFD0EF87C007F03BF7F7ECD9DD561908FFCC7F8000002800;
defparam prom_inst_22.INIT_RAM_0A = 256'hFE21FE000000A00000000C83FFC06600801FE467FFFF89633E0D9AA3FF98FF00;
defparam prom_inst_22.INIT_RAM_0B = 256'hF0F9544FFC43FC000001400000003807FFA00038007FC8CFFEEB703D203830AF;
defparam prom_inst_22.INIT_RAM_0C = 256'hFFFFD36F2773709FF887F800000280000000702FFFA080F200FF919FFFF2EFFA;
defparam prom_inst_22.INIT_RAM_0D = 256'h07F08FFFFF64F5D17CFAA13FF14FF00000058000000AE43FFF00FF8003FE47FF;
defparam prom_inst_22.INIT_RAM_0E = 256'hFD0000001FC13FFFFFF2EAE2B9D5C27FE3DFE000000B00000015C87FFE400000;
defparam prom_inst_22.INIT_RAM_0F = 256'h005701FFFB81F8003F06FFFFFFF059DEF3C1C4FFC7BFC00000160000002B80FF;
defparam prom_inst_22.INIT_RAM_10 = 256'h001C000000AC03FFFC07F8003E6D7FFFBF8E47B0E7A389FF8F7F8000000C0000;
defparam prom_inst_22.INIT_RAM_11 = 256'h3DFE000000380000015805FFF23FF801F19FFFFF7F4A8CDECFA213FF1EFF0000;
defparam prom_inst_22.INIT_RAM_12 = 256'hA6E84FFC63FE00000070000002A00BEFEE7FE007C72FFFFF7F157A779B4427FE;
defparam prom_inst_22.INIT_RAM_13 = 256'hFE5631CE38FA9FF8E7FFC00000F00000074017DF7C3FC00F3EDFFFFCFFB99D2B;
defparam prom_inst_22.INIT_RAM_14 = 256'hC3FFFF637E87215F69DB3FF18FFD400002C000000280279FF80707F879FFFFB1;
defparam prom_inst_22.INIT_RAM_15 = 256'hE0F803FC07FFFEC3E58E613E87203FF63FFEA00001900000C5004FFFE80E0F0F;
defparam prom_inst_22.INIT_RAM_16 = 256'hD0013FFD3FE0000E1FFFFDCE5125CB7CCEAEFFCC7FFF58000320001FCA009E6F;
defparam prom_inst_22.INIT_RAM_17 = 256'h1C007FFF9002FDEC1C0003BE7FFFFB9B66C7CDED9EADFF98FFBED8000E0001FF;
defparam prom_inst_22.INIT_RAM_18 = 256'hE21F78003FFFFFFF2005FF247800001CFFFFF73C0F00BB7B375BFF21FC1F5C00;
defparam prom_inst_22.INIT_RAM_19 = 256'hF29FFD371C1F58006FFFFEE0400BF842F00007F9F7FFEFFD4E53CA78BABFFED3;
defparam prom_inst_22.INIT_RAM_1A = 256'hDFC8EAF7BEDFF2E0C00FD000DFFFFC008017C007E0003DF3EFFFDCC37CB37171;
defparam prom_inst_22.INIT_RAM_1B = 256'h3FFF76371C79F727EFBFE5C30003F8013E3FC001C40DC00FF0001FE79FFFB9B5;
defparam prom_inst_22.INIT_RAM_1C = 256'hC0003F983FFEED82534B9B6FEC3FCB9C000350027CFF000380A1003FE0003FCE;
defparam prom_inst_22.INIT_RAM_1D = 256'h12E001FF80003F307BFDF3706F7E472FCCFFD77000038006DFFC0007026200FF;
defparam prom_inst_22.INIT_RAM_1E = 256'h3F0000061A8007FF00007EE8F3FBE9C7258A723FB1FFACC00601E0001FC0000F;
defparam prom_inst_22.INIT_RAM_1F = 256'h1E02601C7600000C75001FFE0000FDB1E7F7BF80C6BE723E83FF5A038E23200E;
defparam prom_inst_22.INIT_RAM_20 = 256'hDFFD6A171E034008E000001BF0007FFC0001FB67CFEFAEC38EDE7D7C87FEB40D;
defparam prom_inst_22.INIT_RAM_21 = 256'h77727CBC1FFAE64E3F808011C0000035E000FFF80001F6CF9FDDBC54BF39FEFE;
defparam prom_inst_22.INIT_RAM_22 = 256'hFD7FEFC689D9F9F09FF5CEBF3F030041E00000BEF003FFE00005EFBF7F120DF4;
defparam prom_inst_22.INIT_RAM_23 = 256'h0003BF7FFAF6809887B3FBD6FFEB9CDE3E0500C3C000017D4007FFC00009DF3E;
defparam prom_inst_22.INIT_RAM_24 = 256'h003FFE0000075EFFF5EBC071076FFFF4FFD779BC7F0600E780000175A00FFF00;
defparam prom_inst_22.INIT_RAM_25 = 256'h000001F2007FF8000006BCFFEBE6025EB0CFFFF1FFAEF3FC3F8A00ED000002EF;
defparam prom_inst_22.INIT_RAM_26 = 256'hFE10004D0000068000FFF000004D7DFFD3E250A7E5CF7F37FF5DE7FC7F0C006F;
defparam prom_inst_22.INIT_RAM_27 = 256'hFD3753F9FCB8005A00000D4001FFC000009AFBFFA4EA3A1FDFBFFFDFFEBBAFFC;
defparam prom_inst_22.INIT_RAM_28 = 256'hBD57FE1FFB6EB3F9F02000B4000118C003FF800001357FFF48461F2FFF0FF60F;
defparam prom_inst_22.INIT_RAM_29 = 256'hAB91F43F7B3FF67FF6DDE1F1F3D0007800000C0007FF0000046FF3FEDFB34F6F;
defparam prom_inst_22.INIT_RAM_2A = 256'h119BC7EF14D2797EE3DFF47FEDBBC3F1EBA00170000004000FFC000008DFE7FF;
defparam prom_inst_22.INIT_RAM_2B = 256'h3FF0000003B2CFEB7C35777EC7BFE8FFDA7783F3F7A002C0000088001FF80000;
defparam prom_inst_22.INIT_RAM_2C = 256'h00028000FFC0000007458FB892FAFFF7CFFFF3FFA9EF07E7FF0005C000011000;
defparam prom_inst_22.INIT_RAM_2D = 256'hFF80100000050001FF00000006AB9FBDE2FC47EFDDFFE3FF53CB07C7FE400B80;
defparam prom_inst_22.INIT_RAM_2E = 256'h4E2D0FC7BF02C00000080007FE000000074F3EFDCAC6EBBFFCFFC7FEA79607C7;
defparam prom_inst_22.INIT_RAM_2F = 256'hFC799FF28D7B0F8E7E0720000018000FF80000000D9F7FDF09EB577E7CFF8FFD;
defparam prom_inst_22.INIT_RAM_30 = 256'h5CEDDFCDFCF23FE53AF6030C7A0800000520001FF00000001ADE7FFE9F63CF8E;
defparam prom_inst_22.INIT_RAM_31 = 256'h67BCFFFD119F9F9BFFC47FCB75E00F08F41000007F60007FE000000035DCFFFF;
defparam prom_inst_22.INIT_RAM_32 = 256'h000000006B79FFF4CD3F7F37FFC8FF96EFE3970878200003E90000FF80000000;
defparam prom_inst_22.INIT_RAM_33 = 256'h00000FFC0000000059F9FFFD6A51FE7FFE99FF35DFC72E08682800FC018001FF;
defparam prom_inst_22.INIT_RAM_34 = 256'hD080700000001FF8000000005FF1FFFE51B2FCEFFF33FE6FFFCE1E1850400F80;
defparam prom_inst_22.INIT_RAM_35 = 256'hFF9E0E0261BB060010007FE000000000F7F1FFB7537FFFDDFE47FC4FFF8E0E00;
defparam prom_inst_22.INIT_RAM_36 = 256'hFC3FF13D7F1C0C04A141FC0D0000FFC0000000009FE3FFFCD7FFFFB9FC8FF89F;
defparam prom_inst_22.INIT_RAM_37 = 256'h5F3F4FFEF9FFE17A0E381C02429FF07F0001FF8000000001DFE7FF4F77CFBBFF;
defparam prom_inst_22.INIT_RAM_38 = 256'h6FCFFFAD7FFF9FFFF3FFC2F47C781C0E450FC1FD0003FF00000000016FE7FFD4;
defparam prom_inst_22.INIT_RAM_39 = 256'h00000023798FFF9C36F3BFFFE6FF95EC10781C1E067F03F00007FC0000000001;
defparam prom_inst_22.INIT_RAM_3A = 256'h007FE0000000004F778FFF3B69E67FFFDFFF2BCC00F0381D68FC0FE4003FF800;
defparam prom_inst_22.INIT_RAM_3B = 256'hA300FF2000FF80000000001F7B0FFF85B1CC7BFFBFFED7BC01F0381D61807F80;
defparam prom_inst_22.INIT_RAM_3C = 256'h07E03910A601FC4001FE00000000003F3C1FF926E708F7FF7FFDAF7B23E0381C;
defparam prom_inst_22.INIT_RAM_3D = 256'hFFE73B9E4FE47800B4FFF08003FC000000000007CFFFF7EE8E11EEFEBFFA5CF6;
defparam prom_inst_22.INIT_RAM_3E = 256'hB6C7BFFC7FCEF63ECFE83800FFFFE2003FF0000000000039C3FFF9C7FB63DFFE;
defparam prom_inst_22.INIT_RAM_3F = 256'hF8FBC6877BCE7FF8FF9DE87D9FC03001FFFFC0007FE0000000000037E1FFEB16;

pROM prom_inst_23 (
    .DO({prom_inst_23_dout_w[30:0],prom_inst_23_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_23.READ_MODE = 1'b0;
defparam prom_inst_23.BIT_WIDTH = 1;
defparam prom_inst_23.RESET_MODE = "SYNC";
defparam prom_inst_23.INIT_RAM_00 = 256'h0000003FFCFFDAA787DD7FF6FF3B91FF1FD03061FFFF0800FFC000000000003F;
defparam prom_inst_23.INIT_RAM_01 = 256'hFF8000000000007FFCFFCE2B9FD2FFF9FE6C27FF1FC070FFFFFE0001FFC00000;
defparam prom_inst_23.INIT_RAM_02 = 256'hFFF8400FFF0000000000007FF8FD9588BFACFF6BFCD0FF7F3F8019FFFFFC4007;
defparam prom_inst_23.INIT_RAM_03 = 256'h3F8007FFFFE1001FFE000000000001FFF8F7EAD4FDD1FFD7F981FE3F3F803BFF;
defparam prom_inst_23.INIT_RAM_04 = 256'hE685F87E7F00061FFF00003FFC000000000003FFF08FCEC17C23FF8FF303FC3F;
defparam prom_inst_23.INIT_RAM_05 = 256'h0000000000000E7E7700061C3E18007FF800000000003BFFE0531F03EBC4EE9F;
defparam prom_inst_23.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_23.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_24 (
    .DO({prom_inst_24_dout_w[30:0],prom_inst_24_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_24.READ_MODE = 1'b0;
defparam prom_inst_24.BIT_WIDTH = 1;
defparam prom_inst_24.RESET_MODE = "SYNC";
defparam prom_inst_24.INIT_RAM_00 = 256'h000000F7FFFFFFEFE000000003FFE0000000000000000003FFFFFFC0000004EA;
defparam prom_inst_24.INIT_RAM_01 = 256'hFFFFFF00000001FFFFFFFFDFC000000007FF80000000000000000007FFFFFF80;
defparam prom_inst_24.INIT_RAM_02 = 256'h0000003FFFFFFE00000021FFFFFFFFBF800000001FFF0000000000000000001F;
defparam prom_inst_24.INIT_RAM_03 = 256'h000000000000007FFFFFFC0000001D1FFFFFFE7E000000003FFE000000000000;
defparam prom_inst_24.INIT_RAM_04 = 256'hFFF0008000000000000000FFFFFFF80000001C1FFFFFF9FC000000007FF80000;
defparam prom_inst_24.INIT_RAM_05 = 256'h00000003FFE0018000000000000001FFFFFFF8000000181FFFFFF7F000000001;
defparam prom_inst_24.INIT_RAM_06 = 256'hFFFFBF800000000FFFC0030000000000000003FFFFFFF00000001C3FFFFFCFC0;
defparam prom_inst_24.INIT_RAM_07 = 256'h00000A37FFFEFE000000001FFFE7E60000000000000007FFFFFFC00000000C7F;
defparam prom_inst_24.INIT_RAM_08 = 256'hFFFF000000001C1FFFF9FC000000003FFFCFCC000000000000000FFFFFFF8000;
defparam prom_inst_24.INIT_RAM_09 = 256'h0000FFFFFFFE00000000082FFFF7F0000000007FFF9F98001800000000001FFF;
defparam prom_inst_24.INIT_RAM_0A = 256'h7FFF80000003FFFFFFFC00000000081FFFCFC000000001FFFF3F30003C3C0000;
defparam prom_inst_24.INIT_RAM_0B = 256'hFCFCC003FFFF0000010FFFFFFFF800000000083FBFBF8000000003FFFE7E6000;
defparam prom_inst_24.INIT_RAM_0C = 256'h00000FFFF9F9800FFFFE0000063FFFFFFFF000000000097F7EFE0000000007FF;
defparam prom_inst_24.INIT_RAM_0D = 256'hF7F8000000001FFFF3F3003FFFFC00001CFFFFFFFFE0000000000E7FF9FC0000;
defparam prom_inst_24.INIT_RAM_0E = 256'h0000007FDFE0000000003FFFC70383FFFFF80039FFFFFFFFFFE0000000000CFF;
defparam prom_inst_24.INIT_RAM_0F = 256'hFF80000000000CFFBF80000000007FFFCE0F03EFFFC00071FFFFFFFFFFC00000;
defparam prom_inst_24.INIT_RAM_10 = 256'hFFFFFFFFFF00000000100DFEFF0000000000FFFFFC07FFFF9FFC00E1FFFFFFFF;
defparam prom_inst_24.INIT_RAM_11 = 256'h00000381FFFFFFFFFE00000000000DFDFC0000000001FFFFF8070FF83FFC01C1;
defparam prom_inst_24.INIT_RAM_12 = 256'hE0FFC00000000700FFFFFFFFFC00000000000FF7F00000000003FFFFF07FFC00;
defparam prom_inst_24.INIT_RAM_13 = 256'h000FFFFFC0FC300000020E01FFFFFFFFF800000000000DCFE00000000007FFFF;
defparam prom_inst_24.INIT_RAM_14 = 256'h00000000001FFFFF83E3800000041C03FFFFFFFFF000000000000FBF80000000;
defparam prom_inst_24.INIT_RAM_15 = 256'h000019FC00000000003FFFFC3F0000000007FEB7FFFFFFFFC000000000000EFF;
defparam prom_inst_24.INIT_RAM_16 = 256'h8001C000000007F800000000007FFFF7FCF000000010356FFFFFFFFF8000C000;
defparam prom_inst_24.INIT_RAM_17 = 256'hFFFFFFFF0003800000000FE00000000000FFFFFFE7E000000030059FFFFFFFFF;
defparam prom_inst_24.INIT_RAM_18 = 256'h019FEFFFFFFFFFFE0007800000003F800000000001FFFFFF3E00000000F8033F;
defparam prom_inst_24.INIT_RAM_19 = 256'h3800000003FFD3FFFFFFFFFC000F000000001F000000000003FFFFFEFE000000;
defparam prom_inst_24.INIT_RAM_1A = 256'h0FFFFFDDE000000007FFAFFFFFFFFFF8001F000000005C000000000007FFFFF3;
defparam prom_inst_24.INIT_RAM_1B = 256'h000000001FFFFF77F80000000DFBDBFFFFFFFFF0003F00000000580000000000;
defparam prom_inst_24.INIT_RAM_1C = 256'h00002000000004003FFFFDFFF900000007FF9FFFFFFFFFE0007E004000000000;
defparam prom_inst_24.INIT_RAM_1D = 256'h01FE08C0000040000000F8007FFFDE17C00000000FFF3FFFFFFFFFC000FE0860;
defparam prom_inst_24.INIT_RAM_1E = 256'hFFFFFF0003FC08C0000040000001F000FFFF7FA1F0000001FFFF3FFFFFFFFF80;
defparam prom_inst_24.INIT_RAM_1F = 256'hFFFEFFFFFFFFFE0007FC0980000040000007C001FFF9FFE0E0000007FFFE7FFF;
defparam prom_inst_24.INIT_RAM_20 = 256'h0800000FFFFFFFFFFFFFFC000FF819800000C000001F8003FFFFFFF00000000F;
defparam prom_inst_24.INIT_RAM_21 = 256'hFFBFFFFE0000001FFFFFFFFFFFFFF8001FF81B0000008000003F0007FFEFFFF8;
defparam prom_inst_24.INIT_RAM_22 = 256'h038C001FFEFFFFFE0000001FFFFFFFFFFFFFF0003FF01F800000800001E6000F;
defparam prom_inst_24.INIT_RAM_23 = 256'h000100000718003FFFFFFFFE00000077FFFEEFFFFFFFE0007FF01F0002018000;
defparam prom_inst_24.INIT_RAM_24 = 256'hFFE03E00000100001E30007FF7FFFFFF000000EFFFFDFFFFFFFFC000FFF01F00;
defparam prom_inst_24.INIT_RAM_25 = 256'hFFFF0003FFC0190000030000786000FEDFFFFFFF000000FFFFFCFFFFFFFF8001;
defparam prom_inst_24.INIT_RAM_26 = 256'hFFF9FFFFFFFE0007FF80180000020000E0C001FEFFFFFFF38000007FFFFDFFFF;
defparam prom_inst_24.INIT_RAM_27 = 256'hC800003FFFF1FFFFFFFC000FFF00380000020003C18003EBFFFFFFFF800000BF;
defparam prom_inst_24.INIT_RAM_28 = 256'hFFFFF91F0400007FFFF3FFFFFFF8001FFE0030000004000703000F9FFFFFFFFF;
defparam prom_inst_24.INIT_RAM_29 = 256'h1C003F7FFFFFF0C60400007FFFE7FFFFFFF0003FFC0030000004001C0E001F5F;
defparam prom_inst_24.INIT_RAM_2A = 256'h040401E0180079FFFFFFFC2087C000FFFFDFBFFFFFE000FFF800300000040070;
defparam prom_inst_24.INIT_RAM_2B = 256'hE000600000083D007000EBFFFFFFFC10070001FFFF8FFFFFFFC001FFF0002000;
defparam prom_inst_24.INIT_RAM_2C = 256'hFF0007FFC00060000007FD00E001CFFFFFFFFC1003E300FFFFBFFFFFFF8003FF;
defparam prom_inst_24.INIT_RAM_2D = 256'hFEBFFFFFFE000FFF80006000000FDF01C0079FFFFFFFDC2003E401FFFF5FFFFF;
defparam prom_inst_24.INIT_RAM_2E = 256'h03C1E1FFFDFFFFFFFC001FFF00004000007FCE01800EFFFFFFFFF00003C083FF;
defparam prom_inst_24.INIT_RAM_2F = 256'hFFE0300001E1F9FFFB7FFFFFF8003FFE0000C000007FCE83000EFFFFFFFF6000;
defparam prom_inst_24.INIT_RAM_30 = 256'h007FFFFFFFC0100003F8FFFFF6FFFFFFF0007FFC0000C00000FFE686001BFFFF;
defparam prom_inst_24.INIT_RAM_31 = 256'h07FFE31C00DFFFFFEF80000001C4EBFFE5FFFFFFE000FFF80000800203FFE78C;
defparam prom_inst_24.INIT_RAM_32 = 256'h000100000FFFF378007FFCFFBE00000001C1FFFFCFFFFFFFC001FFF000008000;
defparam prom_inst_24.INIT_RAM_33 = 256'h0007FFC0000100001FFFF3B803FFEC3FF000000001D3FFFF9FFFFFFF8003FFE0;
defparam prom_inst_24.INIT_RAM_34 = 256'h2FFFFFFE000FFF80000200001FFFF9C007FFDC3F8001000001FFFFFFBFFFFFFF;
defparam prom_inst_24.INIT_RAM_35 = 256'h00FFFFFC5FFFFFF8001FFF00000200003FFFF8E01FFFFC3C0000000001FBFFFF;
defparam prom_inst_24.INIT_RAM_36 = 256'h0000000000FFFFF8BFFFFFF0003FFE0000060000FFFFFCE039FFC83C00000000;
defparam prom_inst_24.INIT_RAM_37 = 256'h83FF81000000000001FFFFF1FFFFFFE0007FFC0000060001FFFFFD7063FEE208;
defparam prom_inst_24.INIT_RAM_38 = 256'hFFFFFF3C000188040000000001FFFFE37FFFFFC000FFF800000C0001FFFFFF31;
defparam prom_inst_24.INIT_RAM_39 = 256'h000C0003F3FFFF8C010010000000000201EFFF86FFFFFF8001FFF00000070003;
defparam prom_inst_24.INIT_RAM_3A = 256'h07FFC0000018000FC3FFFF84000000000000000201FFFF0DFFFFFF0003FFE000;
defparam prom_inst_24.INIT_RAM_3B = 256'hFFFFFC000FFF80000010000FC7FFDFC2000000000000000601EFF81BFFFFFE00;
defparam prom_inst_24.INIT_RAM_3C = 256'h01FF802FFFFFF8001FFF00000038000C07FF9FE0000000000000000301FFE017;
defparam prom_inst_24.INIT_RAM_3D = 256'h0000000201FF805FFFFFF0003FFE00000030001C07FFFFF00000000000000003;
defparam prom_inst_24.INIT_RAM_3E = 256'h000000000000000731FE00BFFFFFE0007FFC00000030001807FFE7F880000000;
defparam prom_inst_24.INIT_RAM_3F = 256'h0FFFF8FC000000000001000301FC01FFFFFFC000FFF800000060006007FFE3F8;

pROM prom_inst_25 (
    .DO({prom_inst_25_dout_w[30:0],prom_inst_25_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_25.READ_MODE = 1'b0;
defparam prom_inst_25.BIT_WIDTH = 1;
defparam prom_inst_25.RESET_MODE = "SYNC";
defparam prom_inst_25.INIT_RAM_00 = 256'h00C000401FFFF0FE100000000000000381F803FFFFFF8001FFF00000006020E0;
defparam prom_inst_25.INIT_RAM_01 = 256'hFFC00000008001D81FFFE00E10000007C000000311E00FFFFFFF0001FFE00000;
defparam prom_inst_25.INIT_RAM_02 = 256'hFFFC0007FF800000018001BE3FFFFC3E1000000C0FC1000723801FFFFFFE0003;
defparam prom_inst_25.INIT_RAM_03 = 256'h3E00FFFFFFF8000FFF000000018001BE3FFFFE6F80784070FC6000071F007FFF;
defparam prom_inst_25.INIT_RAM_04 = 256'hFC400607FC01FFFFFFF0001FFE0000000300013F3FFFFFEF807F1FC1F8C10703;
defparam prom_inst_25.INIT_RAM_05 = 256'hC201FB8FFC630607FC0FFFFFFFE0003FFC0000000200073F9FFFFFE18046FF80;
defparam prom_inst_25.INIT_RAM_06 = 256'hF3FDF9FBC107FBFE7DC00607F31F7FFFFFC0007FF80000000401033FCFFFFFFE;
defparam prom_inst_25.INIT_RAM_07 = 256'h0800069FF9FB41FF8004FFF7EDA38E0FE73EFFFFFF8000FFF00000000400033F;
defparam prom_inst_25.INIT_RAM_08 = 256'hC00000000900060FFCFC0010990AFF91F8C00E0F847FFFFFFF0001FFE0000000;
defparam prom_inst_25.INIT_RAM_09 = 256'hFC0007FF8000000012000607F6FFE000D917EF8FB0C31E0F0177FFFFFE0003FF;
defparam prom_inst_25.INIT_RAM_0A = 256'h45FFFFFFF8000FFF0000000011000601EF7FC000E927C783B9C00F0E116FFFFF;
defparam prom_inst_25.INIT_RAM_0B = 256'hFC733F1E077FFFFFF0001FFE00000000200002001FBAC08029C7C609DA039F1E;
defparam prom_inst_25.INIT_RAM_0C = 256'hACB7C719EFC5DC1C1EFFFFFFE0003FFC00000000600003002E9D8000CAD76F01;
defparam prom_inst_25.INIT_RAM_0D = 256'hDE460001E416C613FF8786583FFFFFFFC000FFF80000000044000300735F0001;
defparam prom_inst_25.INIT_RAM_0E = 256'h800005837F800001C56D0E31FFE78E3077FFFFFF8001FFF000000000C0000501;
defparam prom_inst_25.INIT_RAM_0F = 256'h000000038000018EFE600001EF981C61DF8F3C50DFFFFFFF0003FFE000000001;
defparam prom_inst_25.INIT_RAM_10 = 256'h000FFF800000001B00000283FDC000004DF794C3FF77DDA7FFFFFFFE0007FFC0;
defparam prom_inst_25.INIT_RAM_11 = 256'hFFFFFFF8001FFF000000003200000207F1E000008BEE09C3FB8F9F0FFFFFFFFC;
defparam prom_inst_25.INIT_RAM_12 = 256'h1FC7FE7BFFFFFFF0003FFE000000006600000456E7F000001FC00E87FEFFBF3D;
defparam prom_inst_25.INIT_RAM_13 = 256'h0F802AF83783F6F7FFFFFFE0007FFC000000004E000008F9CFF800000F801D3E;
defparam prom_inst_25.INIT_RAM_14 = 256'h7FFC00080681A5B072DF3EEFFFFFFFC000FFF800000000CC000010B30FFC0018;
defparam prom_inst_25.INIT_RAM_15 = 256'h0200031CFFF8001046878BC067E7FDFFFFFFFF8001FFF000000000C8010011C6;
defparam prom_inst_25.INIT_RAM_16 = 256'h0000013000000E33FFF0000004025780CFF3FFFFFFFFFF0003FFE00000000190;
defparam prom_inst_25.INIT_RAM_17 = 256'h0FFF80000000002000011867FFF000200406E208B3E3FEFF3FFFFE0007FFC000;
defparam prom_inst_25.INIT_RAM_18 = 256'hFFFFF8001FFF000000000060000230CFFFE000400501C001079FFFFE7FFFFC00;
defparam prom_inst_25.INIT_RAM_19 = 256'h3793AFFFFFFFF0003FFE0000000000C0000461BFFFC00080052F80422F9BD7FF;
defparam prom_inst_25.INIT_RAM_1A = 256'h0DCA6198631B3FFFFFFFE0007FFC0000000000800009877FFF8001008D6730CC;
defparam prom_inst_25.INIT_RAM_1B = 256'hFC0000080918C9C2934FDFFFFFFFC000FFF800000000010000130EFFFE0000A0;
defparam prom_inst_25.INIT_RAM_1C = 256'hC04833FFF80000400E3243C337ADBFFFFFFF8001FFF0000000000100602619FF;
defparam prom_inst_25.INIT_RAM_1D = 256'h0000060080906FFFF00000100A2481E225313FFFFFFF0003FFE0000000000200;
defparam prom_inst_25.INIT_RAM_1E = 256'hFF800000000004011520DFFFC0007CA02A6902866F7C1FFFFFFE0007FFC00000;
defparam prom_inst_25.INIT_RAM_1F = 256'hFFF8001FFF0000000000080064C0CFFF800FFD42185B000CE7239FFFFFFC000F;
defparam prom_inst_25.INIT_RAM_20 = 256'hFF043FFFFFF0003FFE00000000001800C903E707007F8DC6105C081CCE023FFF;
defparam prom_inst_25.INIT_RAM_21 = 256'h41C0C4DF9CF03FFFFFE0007FFC00000000003001920FF80601B808C454B03A0D;
defparam prom_inst_25.INIT_RAM_22 = 256'h1FEDFE943801899FCF003FFFFFC000FFF800000000003003263DF80407F15C8C;
defparam prom_inst_25.INIT_RAM_23 = 256'h983478C039001E9C2807133AE2401FFFFF8001FFF00000000000600A4C3E7838;
defparam prom_inst_25.INIT_RAM_24 = 256'h0000802B30001BC0042006B0801C2A77E3804FFFFF0003FFE00000000000C015;
defparam prom_inst_25.INIT_RAM_25 = 256'h800000000001001660058BC011800F7050F054FBE340DFFFFE0007FFC0000000;
defparam prom_inst_25.INIT_RAM_26 = 256'hF8001FFF000000000003003C40130F81F5B18FE4410089E6E7407FFFFC000FFF;
defparam prom_inst_25.INIT_RAM_27 = 256'hE0967FFFF0003FFE38000000000200788066D703F7BF1FA1A00303C4E2807FFF;
defparam prom_inst_25.INIT_RAM_28 = 256'h80080BFCC1603FFFE0007FFC18000000000400F100CFF60FEEFE7D60800E05DE;
defparam prom_inst_25.INIT_RAM_29 = 256'h083C3C63400035F9E2E19FFFC000FFF800000000000401E2018F6E1E9EED8DB1;
defparam prom_inst_25.INIT_RAM_2A = 256'h1380787801F805418000EBD1FC2087FF8001FFF000000000000803E60901DC3F;
defparam prom_inst_25.INIT_RAM_2B = 256'h00320E183FE0E0D037801D428001D5E370908FFF0007FFE0000000000018070C;
defparam prom_inst_25.INIT_RAM_2C = 256'h0000000000241C307F01C02000002D8280005BCD03F09FFE000FFFC000000000;
defparam prom_inst_25.INIT_RAM_2D = 256'h003BFF018000000000403960F803804000003985000EFD9D93B07FFC001DFFB0;
defparam prom_inst_25.INIT_RAM_2E = 256'hC3FFFFF00077FE03E000000000807241F20F008000007985000FF21FB379FFF8;
defparam prom_inst_25.INIT_RAM_2F = 256'h00F1F83DD209FFE000EFFC07E000000001806483E00E20000000F9C80047EE37;
defparam prom_inst_25.INIT_RAM_30 = 256'h0005F75801AFE06FE2C07F8001CFFA1FE00000000100C90E401C40000000F50A;
defparam prom_inst_25.INIT_RAM_31 = 256'h00F00000000BE3140347802FAE6FFF00039FFE3FC00000000300120FC0780000;
defparam prom_inst_25.INIT_RAM_32 = 256'h0404483801E000000017C220068A00FDCFFFFE00073FFE7F800000000600241C;
defparam prom_inst_25.INIT_RAM_33 = 256'hC60000000888907003C40000000F8FE8053001EBDFFFFC000C7FFFFF02000000;
defparam prom_inst_25.INIT_RAM_34 = 256'h31FFFFFFC4000000111120E0071C0000001F07602E0800C9FDFFF80018FFFFFF;
defparam prom_inst_25.INIT_RAM_35 = 256'hD03DE00063FFFFFF80000000100261E00E3C0000003E0ED0BC301DD5FC7FF000;
defparam prom_inst_25.INIT_RAM_36 = 256'h0DC01CB9D31BE000C7FFFFEF000000002080C1C01C780000007D1EA0246026D9;
defparam prom_inst_25.INIT_RAM_37 = 256'h03FC0D4458802AF7D78F800187FFFFDF100000004101838038F0000000FA0F85;
defparam prom_inst_25.INIT_RAM_38 = 256'hC784000007F82D03F78077FFE9FF00030FFFFFDF0000000042238600E1C20000;
defparam prom_inst_25.INIT_RAM_39 = 256'h088E0C03840C00000FF80BC3ED00EEFFDFFE00061FFFFFFE0000000084470E01;
defparam prom_inst_25.INIT_RAM_3A = 256'h00000003111C1C07081800003FF04E03B6101DBFFFBE000C3FFFFFFE00000001;
defparam prom_inst_25.INIT_RAM_3B = 256'hFFFFFFB8000000020238180E703000007FE080839C961ABFEF7C00187FFFFFDC;
defparam prom_inst_25.INIT_RAM_3C = 256'hFFE00031FFFFFF78000000040070300C7E600000FF809003810EEE3FFFF00030;
defparam prom_inst_25.INIT_RAM_3D = 256'h0C03BE7FFFC00063FFFFFFF00000000900A0300BFE800001FF80A100018DDD7F;
defparam prom_inst_25.INIT_RAM_3E = 256'hFE109DE628AFFE7B7F8000FFFFFFFFE00000001A81406017D9000003FF00C217;
defparam prom_inst_25.INIT_RAM_3F = 256'h0000000FFC2038E6515FE667FF0001FFFFFFFF620000001443C0400318000007;

pROM prom_inst_26 (
    .DO({prom_inst_26_dout_w[30:0],prom_inst_26_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_26.READ_MODE = 1'b0;
defparam prom_inst_26.BIT_WIDTH = 1;
defparam prom_inst_26.RESET_MODE = "SYNC";
defparam prom_inst_26.INIT_RAM_00 = 256'h2F0080F000000017F8499862B0FFCFC3FE0003DFFFFFFEC40000002887808060;
defparam prom_inst_26.INIT_RAM_01 = 256'h000000E21E8100840000000FF081BC25FBFF8FB3FC0007BFFFFFFD8000000071;
defparam prom_inst_26.INIT_RAM_02 = 256'hFFFFFE00000000C03F0001880000001FE2007003D7FF2373F8000F7FFFFFFF00;
defparam prom_inst_26.INIT_RAM_03 = 256'hE0003FFFFFFFFC00000000807E0207300000003F8400746167FA4FF7F0001EFF;
defparam prom_inst_26.INIT_RAM_04 = 256'hAEFD1BF7C0007DFFFFFFF84000000180FC0606600000007F0812E1F0DFFB8FF7;
defparam prom_inst_26.INIT_RAM_05 = 256'h7040EF6BBFF272F78000F787FFFFF8800000034578040300000005FE3062E832;
defparam prom_inst_26.INIT_RAM_06 = 256'hFF0037F8E085EE9FDFC5F4EB8001EE0FFFFFF10000000689F000C00003000BFC;
defparam prom_inst_26.INIT_RAM_07 = 256'hE012FFFFFE00FFF14205DDADBEAE2CEE0003D81FFFFFE20000000117A009F9FF;
defparam prom_inst_26.INIT_RAM_08 = 256'h000004DF4010000FF001FFE28401D86FFD502DEC0007C03FFFFFC4000000022F;
defparam prom_inst_26.INIT_RAM_09 = 256'hFFFF9000000009BE00309007C007FFC40809DCF7EAA1F9C8000F807FFFFFC800;
defparam prom_inst_26.INIT_RAM_0A = 256'h003E01FFFFFF20000000137C00200000801FFB980009A97FD5E37B60001F00FF;
defparam prom_inst_26.INIT_RAM_0B = 256'hEF82F7C0007C03FFFFFE4000000007F800600038007FF730010D90FFE7C5F360;
defparam prom_inst_26.INIT_RAM_0C = 256'h0000575F9984F78000F807FFFFFC800000000FD0006080F200FFEE60000423F7;
defparam prom_inst_26.INIT_RAM_0D = 256'h07FF70000099FDF3231DEF0001F00FFFFFF9800000001BE000C0FF8003FFB800;
defparam prom_inst_26.INIT_RAM_0E = 256'h028000001FFEC000001EFBE6063BDE0003E01FFFFFF30000000037C001C00000;
defparam prom_inst_26.INIT_RAM_0F = 256'h0000FF00048000003FF90000001CFFDE8C3FFC0007C03FFFFFE6000000007F80;
defparam prom_inst_26.INIT_RAM_10 = 256'hFFDC00000003FE00010000003F92800040475FBD187FF8000F807FFFFFEC0000;
defparam prom_inst_26.INIT_RAM_11 = 256'h3E01FFFFFFB800000007FE0008000001FE600000808EBCEF30DFF0001F00FFFF;
defparam prom_inst_26.INIT_RAM_12 = 256'h5B1FC0007C01FFFFFF700000001FFC1012000007F8D0000080FD7B9465BFE000;
defparam prom_inst_26.INIT_RAM_13 = 256'h01E67ED1C71D8000F8043FFFFEF00000003FF8208400000FC120000300799EE8;
defparam prom_inst_26.INIT_RAM_14 = 256'h3C00009C8207BF20966D0001F0033FFFFCC00000007FF860080007FF8600004E;
defparam prom_inst_26.INIT_RAM_15 = 256'h200003FFF800013C198F5D4178760007C0019FFFFD900000C0FFF00018000FF0;
defparam prom_inst_26.INIT_RAM_16 = 256'hC7FFC0034000000FE000023107373B8330F6000F8000C7FFFB20001FC1FFE190;
defparam prom_inst_26.INIT_RAM_17 = 256'hEC007FFF8FFF021BE00003BF800004641EE60C126374001F004047FFF60001FF;
defparam prom_inst_26.INIT_RAM_18 = 256'h1FE0C7FFDFFFFFFF1FFE009B8000001F000008C03FE7BCA4C2A0003E03E0C3FF;
defparam prom_inst_26.INIT_RAM_19 = 256'h0B4001C8FFE0C7FFBFFFFEE03FFC05BD000007FE0800110B7F83D5C7036000EC;
defparam prom_inst_26.INIT_RAM_1A = 256'hDF581F180BC0031FC7F04FFF7FFFFC007FF82FF800003DFC1000232E7FFD4F8E;
defparam prom_inst_26.INIT_RAM_1B = 256'hC00089573FFE3E381780063F0FFC47FEFFFFC000BBF0BFF000001FF86000462D;
defparam prom_inst_26.INIT_RAM_1C = 256'h00003FE7C001115A5CD66BF008000C7C1FFCCFFDFFFF00017FD4FFC000003FF1;
defparam prom_inst_26.INIT_RAM_1D = 256'hED1FFE0000003FCF8402085078E7BFC0300018F03FFC5FFBDFFC0002FD97FF00;
defparam prom_inst_26.INIT_RAM_1E = 256'h3F000001E57FF80000007F1F0C040C07FA278CC0780033C07FFE5FFB1FC00004;
defparam prom_inst_26.INIT_RAM_1F = 256'hFFFD1FEC7600000389FFE0000000FE7E18084A83F9C18DC0B0006603FFFC9FF6;
defparam prom_inst_26.INIT_RAM_20 = 256'h8001981BFFFD3FE8E000000407FF80000001FCF830108EC773218281E000CC0F;
defparam prom_inst_26.INIT_RAM_21 = 256'hA98F030380032077FFFE7FD1C000000A3FFF00000001F9F06020CC5F4CC70101;
defparam prom_inst_26.INIT_RAM_22 = 256'h028327FFF622060C800640CFFFFEFF81E00000403FFC00000005F3C080C151FB;
defparam prom_inst_26.INIT_RAM_23 = 256'h0003CF80050A41FF7844040A000C811FFFFCFF03C0000081FFF800000009E7C1;
defparam prom_inst_26.INIT_RAM_24 = 256'hFFC000000007BF000A1443FEF08800140019023FFFFDFF0780000103FFF00000;
defparam prom_inst_26.INIT_RAM_25 = 256'h0000000FFF80000000077F00141907F54B0000300032047FFFF9FF0D0000020F;
defparam prom_inst_26.INIT_RAM_26 = 256'hFFF7FF8D0000007FFF000000004EFE002C525FF812500060006408FFFFFBFF8F;
defparam prom_inst_26.INIT_RAM_27 = 256'h019063FFFFF7FF9A0000007FFE000000009DFC0058BA26E020A0005000C831FF;
defparam prom_inst_26.INIT_RAM_28 = 256'h43E001000220C7FFFFEFFF34000001FFFC000000013B7800B22C26C001200880;
defparam prom_inst_26.INIT_RAM_29 = 256'h5219FB4086C00A0004410FFFFFCFFF78000027FFF80000000473FC0121317C90;
defparam prom_inst_26.INIT_RAM_2A = 256'h11EBF810F0F246811C200C0008821FFFFF9FFE70000047FFF000000008E7F800;
defparam prom_inst_26.INIT_RAM_2B = 256'hC000000003D2F01B72758C813840180010043FFFFF9FFCC000009FFFE0000000;
defparam prom_inst_26.INIT_RAM_2C = 256'h0002FFFF0000000007A5F07F25FB08083000100034087FFFFF3FF9C000017FFF;
defparam prom_inst_26.INIT_RAM_2D = 256'hFF7FE0000004FFFE00000000076BE0C21AFFB810220020006810FFFFFE3FF380;
defparam prom_inst_26.INIT_RAM_2E = 256'hA043FFFFFEFD0000000FFFF80000000006CFC1023BDF544003004000D021FFFF;
defparam prom_inst_26.INIT_RAM_2F = 256'h038700034187FFFFFDF82000001FFFF0000000000E9F8020EFEDA88183008001;
defparam prom_inst_26.INIT_RAM_30 = 256'h651E6032030E0006830FFFFFF9F00000052FFFE0000000001DDF800093763071;
defparam prom_inst_26.INIT_RAM_31 = 256'h7BBF0001E4784064003C000D061FFFFFF3E000007F5FFF80000000003BDF0002;
defparam prom_inst_26.INIT_RAM_32 = 256'h00000000777E0007B2B080C80038001A081FFFFFF7C00003FF7FFF0000000000;
defparam prom_inst_26.INIT_RAM_33 = 256'hFFFFF0000000000065FE000F957E01800078002C103FFFFFE7C800FFFEFFFE00;
defparam prom_inst_26.INIT_RAM_34 = 256'hCF007FFFFFFFE0000000000067FE0003EDED031000F00058203FFFFFCF800FFF;
defparam prom_inst_26.INIT_RAM_35 = 256'h807FFFFDDE03F9FFFFFF800000000000CFFE0041F380002201E000A0407FFFFF;
defparam prom_inst_26.INIT_RAM_36 = 256'h0280028180FFFFFB9E3603FFDFFF000000000000CFFC0007D600004603C00140;
defparam prom_inst_26.INIT_RAM_37 = 256'h6080B00105800703F1FFFFFD3C680FFFFFFE0000000000018FF8009F58204400;
defparam prom_inst_26.INIT_RAM_38 = 256'h9FF00079800060000B000E07E3FFFFF138E03FFFFFFC0000000000019FF8003E;
defparam prom_inst_26.INIT_RAM_39 = 256'h0000002389F0005FC90C400016001C0FEFFFFFE179A0FFFDFFF8000000000001;
defparam prom_inst_26.INIT_RAM_3A = 256'hFF8000000000004F8FF000AD961980003C00380FFFFFFFE31743FFFBFFC00000;
defparam prom_inst_26.INIT_RAM_3B = 256'h9DFFFFFFFF0000000000001F87F0016A4E3384007800F03FFFFFFFE31EFFFFFF;
defparam prom_inst_26.INIT_RAM_3C = 256'hFFFFFEEF9BFFFFBFFE0000000000003FC3E006B998F70800F001E07CDFFFFFE3;
defparam prom_inst_26.INIT_RAM_3D = 256'h400703E1BFFBFFFF87FFFF7FFC00000000000007F000097331EE1101E003C0F9;
defparam prom_inst_26.INIT_RAM_3E = 256'hCF384003000E07C13FF7FFFFFFFFFFFFC000000000000039FC0005FC479C2001;
defparam prom_inst_26.INIT_RAM_3F = 256'hFF003F739E318006001C0F827FFFFFFFFFFFFBFF8000000000000037FE001FF9;

pROM prom_inst_27 (
    .DO({prom_inst_27_dout_w[30:0],prom_inst_27_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_27.READ_MODE = 1'b0;
defparam prom_inst_27.BIT_WIDTH = 1;
defparam prom_inst_27.RESET_MODE = "SYNC";
defparam prom_inst_27.INIT_RAM_00 = 256'h0000003FFF003DCE5C62800A00385E00FFEFFFFFFFFFF7FF000000000000003F;
defparam prom_inst_27.INIT_RAM_01 = 256'h000000000000007FFF00739CB8CD00040063B800FFFFFFFFFFFFFFFE00000000;
defparam prom_inst_27.INIT_RAM_02 = 256'hFFFF7FF0000000000000007FFF03EE72F193009800CF4080FFFFFFFFFFFFFFF8;
defparam prom_inst_27.INIT_RAM_03 = 256'hFFFFFFFFFFFEFFE000000000000001FFFF0F9565632E003001BE81C0FFFFFFFF;
defparam prom_inst_27.INIT_RAM_04 = 256'h067A0781FFFFFE1FFFFFFFC000000000000003FFFF6A31D6C1DC0060037D03C0;
defparam prom_inst_27.INIT_RAM_05 = 256'h0000000000000F81F7FFFE1C3FFFFF800000000000003BFFFFECE1DD933B1140;
defparam prom_inst_27.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_27.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_28 (
    .DO({prom_inst_28_dout_w[30:0],prom_inst_28_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_28.READ_MODE = 1'b0;
defparam prom_inst_28.BIT_WIDTH = 1;
defparam prom_inst_28.RESET_MODE = "SYNC";
defparam prom_inst_28.INIT_RAM_00 = 256'hFFFFFF080000001FFFFFFFFFFC001FFFFFFFFFFFFFFFFFFC0000003FFFFFFCE3;
defparam prom_inst_28.INIT_RAM_01 = 256'h000000FFFFFFFE000000003FFFFFFFFFF8007FFFFFFFFFFFFFFFFFF80000007F;
defparam prom_inst_28.INIT_RAM_02 = 256'hFFFFFFC0000001FFFFFFDE000000007FFFFFFFFFE000FFFFFFFFFFFFFFFFFFE0;
defparam prom_inst_28.INIT_RAM_03 = 256'hFFFFFFFFFFFFFF80000003FFFFFF82E0000001FFFFFFFFFFC001FFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_04 = 256'h000FFF7FFFFFFFFFFFFFFF00000007FFFFFF03E0000007FFFFFFFFFF8007FFFF;
defparam prom_inst_28.INIT_RAM_05 = 256'hFFFFFFFC001FFE7FFFFFFFFFFFFFFE00000007FFFFFE07E000000FFFFFFFFFFE;
defparam prom_inst_28.INIT_RAM_06 = 256'h00007FFFFFFFFFF0003FFCFFFFFFFFFFFFFFFC0000000FFFFFFC03C000003FFF;
defparam prom_inst_28.INIT_RAM_07 = 256'hFFF005C80001FFFFFFFFFFE0001819FFFFFFFFFFFFFFF80000003FFFFFF80380;
defparam prom_inst_28.INIT_RAM_08 = 256'h0000FFFFFFE003E00007FFFFFFFFFFC0003033FFFFFFFFFFFFFFF00000007FFF;
defparam prom_inst_28.INIT_RAM_09 = 256'hFFFF00000001FFFFFFC007D0000FFFFFFFFFFF80006067FFE7FFFFFFFFFFE000;
defparam prom_inst_28.INIT_RAM_0A = 256'h80007FFFFFFC00000003FFFFFF8007E0003FFFFFFFFFFE0000C0CFFFC3C3FFFF;
defparam prom_inst_28.INIT_RAM_0B = 256'h03033FFC0000FFFFFEF000000007FFFFFF0007C0407FFFFFFFFFFC0001819FFF;
defparam prom_inst_28.INIT_RAM_0C = 256'hFFFFF00006067FF00001FFFFF9C00000000FFFFFFE00068081FFFFFFFFFFF800;
defparam prom_inst_28.INIT_RAM_0D = 256'h0FFFFFFFFFFFE0000C0CFFC00003FFFFE3000000001FFFFFFC00018007FFFFFF;
defparam prom_inst_28.INIT_RAM_0E = 256'hF00007803FFFFFFFFFFFC00038FC7C000007FFC600000000001FFFFFF8000300;
defparam prom_inst_28.INIT_RAM_0F = 256'h007FFFFFE00003007FFFFFFFFFFF800031F0FC10003FFF8E00000000003FFFFF;
defparam prom_inst_28.INIT_RAM_10 = 256'h0000000000FFFFFFC0000201FFFFFFFFFFFF000003F800006003FF1E00000000;
defparam prom_inst_28.INIT_RAM_11 = 256'hFFFFFC7E0000000001FFFFFF80000203FFFFFFFFFFFE000007F8F007C003FE3E;
defparam prom_inst_28.INIT_RAM_12 = 256'h1F003FFFFFFFF8FF0000000003FFFFFF0000000FFFFFFFFFFFFC00000F8003FF;
defparam prom_inst_28.INIT_RAM_13 = 256'hFFF000003F03FFFFFFFDF1FE0000000007FFFFFE0000023FFFFFFFFFFFF80000;
defparam prom_inst_28.INIT_RAM_14 = 256'hFFFFFFFFFFE000007C1FFFFFFFFBE3FC000000000FFFFFFC0000007FFFFFFFFF;
defparam prom_inst_28.INIT_RAM_15 = 256'h000007FFFFFFFFFFFFC00003C0FFFFFFFFF80148000000003FFFFFF8000001FF;
defparam prom_inst_28.INIT_RAM_16 = 256'h7FFE3FE000000FFFFFFFFFFFFF80000803FFFFFFFFEFCA90000000007FFF3FF0;
defparam prom_inst_28.INIT_RAM_17 = 256'h00000000FFFC7FC000001FFFFFFFFFFFFF0000001FFFFFFFFFCFFA6000000000;
defparam prom_inst_28.INIT_RAM_18 = 256'hFE60100000000001FFF87F8000001FFFFFFFFFFFFE000000FFFFFFFFFF07FCC0;
defparam prom_inst_28.INIT_RAM_19 = 256'hFFFFFFFFFC002C0000000003FFF0FF0000003FFFFFFFFFFFFC000001FFFFFFFF;
defparam prom_inst_28.INIT_RAM_1A = 256'hF000003FFFFFFFFFF800500000000007FFE0FE0000003FFFFFFFFFFFF800000F;
defparam prom_inst_28.INIT_RAM_1B = 256'hFFFFFFFFE00000FFFFFFFFFFF20424000000000FFFC0FC0000003FFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_1C = 256'h00001FFFFFFFFBFFC00003FFFFFFFFFFF80060000000001FFF81F80000003FFF;
defparam prom_inst_28.INIT_RAM_1D = 256'hFE01F00000003FFFFFFF07FF80003FFFFFFFFFFFF000C0000000003FFF01F000;
defparam prom_inst_28.INIT_RAM_1E = 256'h000000FFFC03F00000003FFFFFFE0FFF0000FFFFFFFFFFFE0000C0000000007F;
defparam prom_inst_28.INIT_RAM_1F = 256'h00010000000001FFF803F00000003FFFFFF83FFE0003FFFFFFFFFFF800018000;
defparam prom_inst_28.INIT_RAM_20 = 256'hFFFFFFF000000000000003FFF007E00000003FFFFFE07FFC0007FFFFFFFFFFF0;
defparam prom_inst_28.INIT_RAM_21 = 256'h007FFFFFFFFFFFE000000000000007FFE007E00000007FFFFFC0FFF8001FFFFF;
defparam prom_inst_28.INIT_RAM_22 = 256'hFC03FFE001FFFFFFFFFFFFE00000000000000FFFC00FE00000007FFFFE01FFF0;
defparam prom_inst_28.INIT_RAM_23 = 256'h0000FFFFF807FFC003FFFFFFFFFFFF880001100000001FFF800FE00000007FFF;
defparam prom_inst_28.INIT_RAM_24 = 256'h001FC0000000FFFFE00FFF800FFFFFFFFFFFFF100002000000003FFF000FE000;
defparam prom_inst_28.INIT_RAM_25 = 256'h0000FFFC003FE0000000FFFF801FFF003FFFFFFFFFFFFF000003000000007FFE;
defparam prom_inst_28.INIT_RAM_26 = 256'h000600000001FFF8007FE0000001FFFF003FFE01FFFFFFFFFFFFFF8000020000;
defparam prom_inst_28.INIT_RAM_27 = 256'hF7FFFFC0000E00000003FFF000FFC0000001FFFC007FFC07FFFFFFFFFFFFFF40;
defparam prom_inst_28.INIT_RAM_28 = 256'hFFFFFFFFFBFFFF80000C00000007FFE001FFC0000003FFF800FFF00FFFFFFFFF;
defparam prom_inst_28.INIT_RAM_29 = 256'h03FFC0FFFFFFFFFFFBFFFF8000180000000FFFC003FFC0000003FFE001FFE03F;
defparam prom_inst_28.INIT_RAM_2A = 256'h0003FE0007FF83FFFFFFFFFFF83FFF0000304000001FFF0007FFC0000003FF80;
defparam prom_inst_28.INIT_RAM_2B = 256'h1FFF80000007FE000FFF07FFFFFFFFFFF8FFFE0000700000003FFE000FFFC000;
defparam prom_inst_28.INIT_RAM_2C = 256'h00FFF8003FFF8000000FFE001FFE1FFFFFFFFFFFFC1CFF0000600000007FFC00;
defparam prom_inst_28.INIT_RAM_2D = 256'h01C0000001FFF0007FFF8000001FFE003FF83FFFFFFFFFFFFC1BFE0000E00000;
defparam prom_inst_28.INIT_RAM_2E = 256'hFC3E1E000380000003FFE000FFFF8000003FFF007FF07FFFFFFFFFFFFC3F7C00;
defparam prom_inst_28.INIT_RAM_2F = 256'hFFFFFFFFFE1E06000780000007FFC001FFFF000000FFFF00FFF1FFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_30 = 256'hFF8FFFFFFFFFFFFFFC0700000F0000000FFF8003FFFF000001FFFF01FFE7FFFF;
defparam prom_inst_28.INIT_RAM_31 = 256'h07FFFF83FF3FFFFFFFFFFFFFFE3B14001E0000001FFF0007FFFF000003FFFF03;
defparam prom_inst_28.INIT_RAM_32 = 256'hFFFE00000FFFFF87FFFFFFFFFFFFFFFFFE3E00003C0000003FFE000FFFFF0000;
defparam prom_inst_28.INIT_RAM_33 = 256'hFFF8003FFFFE00001FFFFFC7FFFFFFFFFFFFFFFFFE2C0000780000007FFC001F;
defparam prom_inst_28.INIT_RAM_34 = 256'hF0000001FFF0007FFFFC00003FFFFFFFFFFFFFFFFFFFFFFFFE00000070000000;
defparam prom_inst_28.INIT_RAM_35 = 256'hFF000003E0000007FFE000FFFFFC00007FFFFFFFFFFFFFFFFFFFFFFFFE040000;
defparam prom_inst_28.INIT_RAM_36 = 256'hFFFFFFFFFF000007C000000FFFC001FFFFF800007FFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFE00000F8000001FFF8003FFFFF80000FFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFE00001F8000003FFF0007FFFFF00001FFFFFFFF;
defparam prom_inst_28.INIT_RAM_39 = 256'hFFF00007FFFFFFFFFFFFFFFFFFFFFFFDFE10007F0000007FFE000FFFFFF80003;
defparam prom_inst_28.INIT_RAM_3A = 256'hF8003FFFFFE00007FFFFFFFFFFFFFFFFFFFFFFFDFE0000FE000000FFFC001FFF;
defparam prom_inst_28.INIT_RAM_3B = 256'h000003FFF0007FFFFFE0000FFFFFFFFFFFFFFFFFFFFFFFF9FE1007FC000001FF;
defparam prom_inst_28.INIT_RAM_3C = 256'hFE007FF0000007FFE000FFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFCFE001FF8;
defparam prom_inst_28.INIT_RAM_3D = 256'hFFFFFFFDFE007FE000000FFFC001FFFFFFC0001FFFFFFFFFFFFFFFFFFFFFFFFC;
defparam prom_inst_28.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFF8CE01FFC000001FFF8003FFFFFFC0003FFFFFFFFFFFFFFFFF;
defparam prom_inst_28.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFEFFFCFE03FF8000003FFF0007FFFFFF80003FFFFFFFFF;

pROM prom_inst_29 (
    .DO({prom_inst_29_dout_w[30:0],prom_inst_29_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_29.READ_MODE = 1'b0;
defparam prom_inst_29.BIT_WIDTH = 1;
defparam prom_inst_29.RESET_MODE = "SYNC";
defparam prom_inst_29.INIT_RAM_00 = 256'hFF0000FFFFFFFFFFFFFFFFFFFFFFFFFC7E07FF0000007FFE000FFFFFFF80007F;
defparam prom_inst_29.INIT_RAM_01 = 256'h003FFFFFFF0000E7FFFFFFFFFFFFFFF83FFFFFFCEE1FFE000000FFFE001FFFFF;
defparam prom_inst_29.INIT_RAM_02 = 256'h0003FFF8007FFFFFFE0001C1FFFFFFFFFFFFFFF3F03EFFF8DC7FFC000001FFFC;
defparam prom_inst_29.INIT_RAM_03 = 256'hC1FFF0000007FFF000FFFFFFFE0003C1FFFFFFFFFF87BF8F039FFFF8E0FFF800;
defparam prom_inst_29.INIT_RAM_04 = 256'h03BFF9F803FFE000000FFFE001FFFFFFFC0003C0FFFFFFFFFF00E03E073EF8FC;
defparam prom_inst_29.INIT_RAM_05 = 256'hFC000070039CF9F803FFC000001FFFC003FFFFFFFC0003C07FFFFFFFFE00007C;
defparam prom_inst_29.INIT_RAM_06 = 256'h0FFFFFFFFE000001823FF9F80CFF8000003FFF8007FFFFFFF80007C03FFFFFFF;
defparam prom_inst_29.INIT_RAM_07 = 256'hF00003E007FFFFFFFE000000125C71F018FF0000007FFF000FFFFFFFF80007C0;
defparam prom_inst_29.INIT_RAM_08 = 256'h3FFFFFFFF00003F003FFFFFFE6000000073FF1F07BFC000000FFFE001FFFFFFF;
defparam prom_inst_29.INIT_RAM_09 = 256'h03FFF8007FFFFFFFE00003F809FFFFFFE60000000F3CE1F0FFF8000001FFFC00;
defparam prom_inst_29.INIT_RAM_0A = 256'hBFC0000007FFF000FFFFFFFFE00003FE10FFFFFFF6000000063FF0F1EFF00000;
defparam prom_inst_29.INIT_RAM_0B = 256'h038CC0E1FF8000000FFFE001FFFFFFFFC00007FFE07FFFFFF600010005FC60E1;
defparam prom_inst_29.INIT_RAM_0C = 256'hF3000000003A23E3FF0000001FFFC003FFFFFFFF800007FFD07FFFFFF7008000;
defparam prom_inst_29.INIT_RAM_0D = 256'h203FFFFFFB200000007879A7FC0000003FFF0007FFFFFFFF800007FF883FFFFF;
defparam prom_inst_29.INIT_RAM_0E = 256'h000003FC807FFFFFFA000000001871CFF80000007FFE000FFFFFFFFF000003FE;
defparam prom_inst_29.INIT_RAM_0F = 256'hFFFFFFFC000003F101FFFFFFF04000000070C3AFE0000000FFFC001FFFFFFFFE;
defparam prom_inst_29.INIT_RAM_10 = 256'hFFF0007FFFFFFFE4000001FC03FFFFFFF20000000088225F80000001FFF8003F;
defparam prom_inst_29.INIT_RAM_11 = 256'h00000007FFE000FFFFFFFFCC000001F80FFFFFFFF4000000007060FF00000003;
defparam prom_inst_29.INIT_RAM_12 = 256'h003801FC0000000FFFC001FFFFFFFF98000003A01FFFFFFFE0000000010040FE;
defparam prom_inst_29.INIT_RAM_13 = 256'hF0001000007C09F80000001FFF8003FFFFFFFFB0000007003FFFFFFFF0000000;
defparam prom_inst_29.INIT_RAM_14 = 256'hFFFFFFFFF90040000120C1F00000003FFF0007FFFFFFFF3000000F00FFFFFFFF;
defparam prom_inst_29.INIT_RAM_15 = 256'h00003C03FFFFFFFFB9000000001803C00000007FFE000FFFFFFFFF3000000E01;
defparam prom_inst_29.INIT_RAM_16 = 256'hFFFFFEC00000700FFFFFFFFFFB010000000C0380000000FFFC001FFFFFFFFE60;
defparam prom_inst_29.INIT_RAM_17 = 256'hF0007FFFFFFFFFC00000E01FFFFFFFFFFB000000001C0700C00001FFF8003FFF;
defparam prom_inst_29.INIT_RAM_18 = 256'h000007FFE000FFFFFFFFFF800001C03FFFFFFFFFFA08000000600C01800003FF;
defparam prom_inst_29.INIT_RAM_19 = 256'h006C700000000FFFC001FFFFFFFFFF000003807FFFFFFFFFFA10000000643800;
defparam prom_inst_29.INIT_RAM_1A = 256'hF200000000E4C00000001FFF8003FFFFFFFFFF00000600FFFFFFFFFFF2000000;
defparam prom_inst_29.INIT_RAM_1B = 256'hFFFFFFFFF600000000B0200000003FFF0007FFFFFFFFFE00000C01FFFFFFFFDF;
defparam prom_inst_29.INIT_RAM_1C = 256'h00300FFFFFFFFFFFF00000000052400000007FFE000FFFFFFFFFFE00001807FF;
defparam prom_inst_29.INIT_RAM_1D = 256'hFFFFF80000601FFFFFFFFFFFF400000002CEC0000000FFFC001FFFFFFFFFFC00;
defparam prom_inst_29.INIT_RAM_1E = 256'h007FFFFFFFFFF80000C03FFFFFFF83FFF40000000081E0000001FFF8003FFFFF;
defparam prom_inst_29.INIT_RAM_1F = 256'h0007FFE000FFFFFFFFFFF00003003FFFFFF003FFE400000000C0E0000003FFF0;
defparam prom_inst_29.INIT_RAM_20 = 256'h0083C000000FFFC001FFFFFFFFFFE00006001FFFFF8073FFEC00000001C1C000;
defparam prom_inst_29.INIT_RAM_21 = 256'hF8000000030FC000001FFF8003FFFFFFFFFFC0000C0007FFFE07F7FFE8000020;
defparam prom_inst_29.INIT_RAM_22 = 256'hE00001FFC000000000FFC000003FFF0007FFFFFFFFFFC000180207FFF80EA3FF;
defparam prom_inst_29.INIT_RAM_23 = 256'h600007FFC60001FFD000000101BFE000007FFE000FFFFFFFFFFF8000300007FF;
defparam prom_inst_29.INIT_RAM_24 = 256'hFFFF0000C00007FFF80001FFF0000000007FF00000FFFC001FFFFFFFFFFF0000;
defparam prom_inst_29.INIT_RAM_25 = 256'h7FFFFFFFFFFE0001800207FFE06001FFA000000000BFE00001FFF8003FFFFFFF;
defparam prom_inst_29.INIT_RAM_26 = 256'h07FFE000FFFFFFFFFFFC0003000C07FE03C001FFA000000000BFC00003FFF000;
defparam prom_inst_29.INIT_RAM_27 = 256'h007900000FFFC001C7FFFFFFFFFC000600180FFC0F0001FF40000000017F8000;
defparam prom_inst_29.INIT_RAM_28 = 256'h4000040000FE00001FFF8003E7FFFFFFFFF8000C00300FF01F0003FF40000200;
defparam prom_inst_29.INIT_RAM_29 = 256'hFFC3C3FE80000A00007E00003FFF0007FFFFFFFFFFF8001800709FE17F1073FE;
defparam prom_inst_29.INIT_RAM_2A = 256'h007FFF87FE07FBFE00001400007F08007FFE000FFFFFFFFFFFF0003000FE3FC0;
defparam prom_inst_29.INIT_RAM_2B = 256'hFFC001C0001FFF2FC87FE3FD00002800006F1000FFF8001FFFFFFFFFFFE000E0;
defparam prom_inst_29.INIT_RAM_2C = 256'hFFFFFFFFFFC0038000FFFFDFFFFFD3FD0001A002C00F6001FFF0003FFFFFFFFF;
defparam prom_inst_29.INIT_RAM_2D = 256'hFFC000FFFFFFFFFFFF80060007FFFFBFFFFFC3FA00010002000F8003FFE0007F;
defparam prom_inst_29.INIT_RAM_2E = 256'h0000000FFF8001FFFFFFFFFFFF000C000DFFFF7FFFFF83FA0000000000060007;
defparam prom_inst_29.INIT_RAM_2F = 256'h000E000201F6001FFF0003FFFFFFFFFFFE0018001FFFDFFFFFFF03F600080000;
defparam prom_inst_29.INIT_RAM_30 = 256'hFFFA03E400400010003F807FFE0007FFFFFFFFFFFE003001BFFFBFFFFFFF03F4;
defparam prom_inst_29.INIT_RAM_31 = 256'hFFFFFFFFFFF407E800800010001000FFFC000FFFFFFFFFFFFC00E0003FFFFFFF;
defparam prom_inst_29.INIT_RAM_32 = 256'hF8038007FFFFFFFFFFE807D801000000000001FFF8001FFFFFFFFFFFF801C003;
defparam prom_inst_29.INIT_RAM_33 = 256'hF9FFFFFFF007000FFFFBFFFFFFF007900A000010000003FFF0003FFFFDFFFFFF;
defparam prom_inst_29.INIT_RAM_34 = 256'hC000FFFFFBFFFFFFE00E001FFFE3FFFFFFE00F9010000020020007FFE0007FFF;
defparam prom_inst_29.INIT_RAM_35 = 256'h21C21FFF8001FFFFFFFFFFFFE03C001FFFC3FFFFFFC00F204000000003800FFF;
defparam prom_inst_29.INIT_RAM_36 = 256'h7000030020E41FFF0003FFFFFFFFFFFFC078003FFF87FFFFFF800F4198000100;
defparam prom_inst_29.INIT_RAM_37 = 256'hFC001E80E100150020707FFE0007FFFFEFFFFFFF80F0007FFF0FFFFFFF001E42;
defparam prom_inst_29.INIT_RAM_38 = 256'hF87BFFFFF8001E80080008000600FFFC000FFFFFFFFFFFFF81C001FFFE3DFFFF;
defparam prom_inst_29.INIT_RAM_39 = 256'h070003FFFBF3FFFFF0003C00100010000001FFF8001FFFFFFFFFFFFF038001FF;
defparam prom_inst_29.INIT_RAM_3A = 256'hFFFFFFFC0E0003FFF7E7FFFFC0003180480160000041FFF0003FFFFFFFFFFFFE;
defparam prom_inst_29.INIT_RAM_3B = 256'h00FFFFFFFFFFFFFC3C0007FF8FCFFFFF80007F000000C1001083FFE0007FFFFF;
defparam prom_inst_29.INIT_RAM_3C = 256'h001FFFC001FFFFFFFFFFFFF878000FFF819FFFFF00007F0000010100000FFFC0;
defparam prom_inst_29.INIT_RAM_3D = 256'h002C0000003FFF8003FFFFFFFFFFFFF0F0000FFC017FFFFE00007E0300120200;
defparam prom_inst_29.INIT_RAM_3E = 256'h0000620010500000807FFF0007FFFFFFFFFFFFE160001FF826FFFFFC00007C00;
defparam prom_inst_29.INIT_RAM_3F = 256'hFFFFFFF00000C70020A0000000FFFE000FFFFFFDFFFFFFE380003FFCE7FFFFF8;

pROM prom_inst_30 (
    .DO({prom_inst_30_dout_w[30:0],prom_inst_30_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_30.READ_MODE = 1'b0;
defparam prom_inst_30.BIT_WIDTH = 1;
defparam prom_inst_30.RESET_MODE = "SYNC";
defparam prom_inst_30.INIT_RAM_00 = 256'h00007FFFFFFFFFE80000E7804300000C01FFFC001FFFFFFBFFFFFFC700007FFF;
defparam prom_inst_30.INIT_RAM_01 = 256'hFFFFFF1C0000FFFFFFFFFFF00000C7C00400000C03FFF8003FFFFFFFFFFFFF8E;
defparam prom_inst_30.INIT_RAM_02 = 256'hFFFFFFFFFFFFFF380001FFFFFFFFFFE000018FC00800040C07FFF0007FFFFFFF;
defparam prom_inst_30.INIT_RAM_03 = 256'h1FFFC001FFFFFFFFFFFFFF700001FFFFFFFFFFC000018F80980000080FFFE000;
defparam prom_inst_30.INIT_RAM_04 = 256'h400000083FFF8003FFFFFFBFFFFFFE600001FFFFFFFFFF8000011E0120000008;
defparam prom_inst_30.INIT_RAM_05 = 256'h00031F84000001087FFF0007FFFFFF7FFFFFFC800003FFFFFFFFFA0000011FC1;
defparam prom_inst_30.INIT_RAM_06 = 256'h00FFC80000021F60000003107FFE000FFFFFFEFFFFFFF90000073FFFFCFFF400;
defparam prom_inst_30.INIT_RAM_07 = 256'h000D000001FF000000023E4201000311FFFC001FFFFFFDFFFFFFFE0000060600;
defparam prom_inst_30.INIT_RAM_08 = 256'hFFFFF800000FFFF00FFE000000063F8002000213FFF8003FFFFFFBFFFFFFFC00;
defparam prom_inst_30.INIT_RAM_09 = 256'hFFFFEFFFFFFFF000000F7FF83FF800000006330004000637FFF0007FFFFFF7FF;
defparam prom_inst_30.INIT_RAM_0A = 256'hFFC001FFFFFFDFFFFFFFE000001FFFFF7FE00000000676800800041FFFE000FF;
defparam prom_inst_30.INIT_RAM_0B = 256'h1004083FFF8003FFFFFFBFFFFFFFC000001FFFC7FF80000000066F0018020C1F;
defparam prom_inst_30.INIT_RAM_0C = 256'h000FA8806008087FFF0007FFFFFF7FFFFFFF8000001F7F0DFF000000000FDC00;
defparam prom_inst_30.INIT_RAM_0D = 256'hF8000000000F020CC00010FFFE000FFFFFFE7FFFFFFF0000003F007FFC000000;
defparam prom_inst_30.INIT_RAM_0E = 256'h007FFFFFE0000000000F0419C00021FFFC001FFFFFFCFFFFFFFE0000003FFFFF;
defparam prom_inst_30.INIT_RAM_0F = 256'hFFF80000007FFFFFC0000000000F0021000003FFF8003FFFFFF9FFFFFFFC0000;
defparam prom_inst_30.INIT_RAM_10 = 256'hFFE3FFFFFFF0000000FFFFFFC00000000018A042000007FFF0007FFFFFF3FFFF;
defparam prom_inst_30.INIT_RAM_11 = 256'hC001FFFFFFC7FFFFFFE0000001FFFFFE000000000031430000000FFFE000FFFF;
defparam prom_inst_30.INIT_RAM_12 = 256'h00003FFF8003FFFFFF8FFFFFFFC0000001FFFFF8000000000002840800001FFF;
defparam prom_inst_30.INIT_RAM_13 = 256'h0019802000007FFF0003FFFFFF0FFFFFFF80000003FFFFF00000000000066010;
defparam prom_inst_30.INIT_RAM_14 = 256'h0000000001F840C00010FFFE0000FFFFFF3FFFFFFF00000007FFF80000000000;
defparam prom_inst_30.INIT_RAM_15 = 256'h1FFFFC0000000000067082800099FFF800007FFFFE6FFFFF3E00000007FFF000;
defparam prom_inst_30.INIT_RAM_16 = 256'h38000000FFFFFFF00000000038C804000119FFF000003FFFFCDFFFE03C000000;
defparam prom_inst_30.INIT_RAM_17 = 256'hF3FF800070000007FFFFFC4000000000E1183200001BFFE000003FFFF9FFFE00;
defparam prom_inst_30.INIT_RAM_18 = 256'h00003FFFE0000000E000007FFFFFFFE000000003C0184000001FFFC000003FFF;
defparam prom_inst_30.INIT_RAM_19 = 256'h043FFE0000003FFFC000011FC00003FFFFFFF80000000004803C2000041FFF00;
defparam prom_inst_30.INIT_RAM_1A = 256'h20270000043FFC0038003FFF800003FF80001FFFFFFFC2000000001180008000;
defparam prom_inst_30.INIT_RAM_1B = 256'h00000088C0000000087FF800F0003FFF00003FFF00007FFFFFFFE00000000042;
defparam prom_inst_30.INIT_RAM_1C = 256'hFFFFC00000000225A020040017FFF003E0003FFE0000FFFE0003FFFFFFFFC000;
defparam prom_inst_30.INIT_RAM_1D = 256'h003FFFFFFFFFC0000000048F800000000FFFE00FC0003FFC2003FFFC000FFFFF;
defparam prom_inst_30.INIT_RAM_1E = 256'hC0FFFFF800FFFFFFFFFF800000001338004000000FFFC03F80003FFCE03FFFF8;
defparam prom_inst_30.INIT_RAM_1F = 256'h0000FFF389FFFFF003FFFFFFFFFF00000000247C000000005FFF81FC00007FF9;
defparam prom_inst_30.INIT_RAM_20 = 256'h7FFE07E00000FFF71FFFFFE00FFFFFFFFFFE000000005138000000003FFF03F0;
defparam prom_inst_30.INIT_RAM_21 = 256'h00000000FFFC1F800001FFEE3FFFFFC01FFFFFFFFFFE0000000123A000000000;
defparam prom_inst_30.INIT_RAM_22 = 256'h00041800000400037FF83F000001FFFE1FFFFF807FFFFFFFFFFA000000028E00;
defparam prom_inst_30.INIT_RAM_23 = 256'hFFFC0000000C3E0000080005FFF07E000003FFFC3FFFFF00FFFFFFFFFFF60000;
defparam prom_inst_30.INIT_RAM_24 = 256'hFFFFFFFFFFF8000000183C000010000BFFE0FC000003FFF87FFFFE03FFFFFFFF;
defparam prom_inst_30.INIT_RAM_25 = 256'hFFFFFC1FFFFFFFFFFFF800000030F8000030000FFFC1F8000007FFF2FFFFFC07;
defparam prom_inst_30.INIT_RAM_26 = 256'h000FFFF2FFFFF83FFFFFFFFFFFB000000021A0000020001FFF83F0000007FFF0;
defparam prom_inst_30.INIT_RAM_27 = 256'hFE0F8000000FFFE5FFFFF0FFFFFFFFFFFF6000000145C1000040002FFF07C000;
defparam prom_inst_30.INIT_RAM_28 = 256'h000000FFFC1F0000001FFFCBFFFFE1FFFFFFFFFFFEC0800003D3C00000C0007F;
defparam prom_inst_30.INIT_RAM_29 = 256'h01E60000000001FFF83E0000003FFF87FFFFC3FFFFFFFFFFFB80000000CE8000;
defparam prom_inst_30.INIT_RAM_2A = 256'hEE0400000F0D8000000003FFF07C0000007FFF8FFFFF8FFFFFFFFFFFF7000000;
defparam prom_inst_30.INIT_RAM_2B = 256'hFFFFFFFFFC0D0004800A0000000007FFE1F80000007FFF3FFFFF1FFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_2C = 256'hFFFC7FFFFFFFFFFFF81A00000004000000000FFFC3F0000000FFFE3FFFFE3FFF;
defparam prom_inst_30.INIT_RAM_2D = 256'h00FFFFFFFFF9FFFFFFFFFFFFF81400000100000000001FFF87E0000001FFFC7F;
defparam prom_inst_30.INIT_RAM_2E = 256'h1F80000001FFFFFFFFF3FFFFFFFFFFFFF83000000420000000003FFF0FC00000;
defparam prom_inst_30.INIT_RAM_2F = 256'h0000FFFC3E00000003FFDFFFFFE7FFFFFFFFFFFFF06000001010000000007FFE;
defparam prom_inst_30.INIT_RAM_30 = 256'h820000000001FFF87C00000007FFFFFFFADFFFFFFFFFFFFFE020000160800000;
defparam prom_inst_30.INIT_RAM_31 = 256'h80400002080000000003FFF0F80000000FFFFFFF80BFFFFFFFFFFFFFC0200001;
defparam prom_inst_30.INIT_RAM_32 = 256'hFFFFFFFF80800000004000000007FFE1F00000000FFFFFFC00FFFFFFFFFFFFFF;
defparam prom_inst_30.INIT_RAM_33 = 256'h03FFFFFFFFFFFFFF82000000008000000007FFC3E00000001FF7FF0001FFFFFF;
defparam prom_inst_30.INIT_RAM_34 = 256'h3FFF800007FFFFFFFFFFFFFF8000000002000000000FFF87C00000003FFFF000;
defparam prom_inst_30.INIT_RAM_35 = 256'h000000003FFC00000FFFFFFFFFFFFFFF000000000C000000001FFF1F80000000;
defparam prom_inst_30.INIT_RAM_36 = 256'h017FFC7E000000007FF800003FFFFFFFFFFFFFFF0000000028000000003FFE3F;
defparam prom_inst_30.INIT_RAM_37 = 256'h80000000027FF8FC00000000FFF000007FFFFFFFFFFFFFFE00000000A0000000;
defparam prom_inst_30.INIT_RAM_38 = 256'h000000060000000004FFF1F800000000FFF00000FFFFFFFFFFFFFFFE00000001;
defparam prom_inst_30.INIT_RAM_39 = 256'hFFFFFFDC060000200000000009FFE3F000000000FFC00003FFFFFFFFFFFFFFFE;
defparam prom_inst_30.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFB0000000400000000003FFC7F000000000FF800007FFFFFFFF;
defparam prom_inst_30.INIT_RAM_3B = 256'h7E00001FFFFFFFFFFFFFFFE0000000100000000007FF0FC000000000FF00000F;
defparam prom_inst_30.INIT_RAM_3C = 256'h000000007C00007FFFFFFFFFFFFFFFC000000040000000000FFE1F8000000000;
defparam prom_inst_30.INIT_RAM_3D = 256'h3FF8FC0000000000780000FFFFFFFFFFFFFFFFF800000080000000001FFC3F00;
defparam prom_inst_30.INIT_RAM_3E = 256'h00000000FFF1F80000000000000001FFFFFFFFFFFFFFFFC60000020000000000;
defparam prom_inst_30.INIT_RAM_3F = 256'h0000000000000001FFE3F00000000000000007FFFFFFFFFFFFFFFFC800000000;

pROM prom_inst_31 (
    .DO({prom_inst_31_dout_w[30:0],prom_inst_31_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_31.READ_MODE = 1'b0;
defparam prom_inst_31.BIT_WIDTH = 1;
defparam prom_inst_31.RESET_MODE = "SYNC";
defparam prom_inst_31.INIT_RAM_00 = 256'hFFFFFFC00000000020000001FFC7E0000000000000000FFFFFFFFFFFFFFFFFC0;
defparam prom_inst_31.INIT_RAM_01 = 256'hFFFFFFFFFFFFFF800000000040000003FF9FC0000000000000001FFFFFFFFFFF;
defparam prom_inst_31.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFFFFF800000000100000007FF3F80000000000000003FFF;
defparam prom_inst_31.INIT_RAM_03 = 256'h000000000001FFFFFFFFFFFFFFFFFE00000000020000000FFE7F000000000000;
defparam prom_inst_31.INIT_RAM_04 = 256'hF9FC0000000001E00003FFFFFFFFFFFFFFFFFC00001000080200001FFCFE0000;
defparam prom_inst_31.INIT_RAM_05 = 256'h0000000000000000080001E3C007FFFFFFFFFFFFFFFFC400000000200400003F;
defparam prom_inst_31.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_31.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[15]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_1)
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(prom_inst_2_dout[0]),
  .I1(prom_inst_3_dout[0]),
  .S0(dff_q_1)
);
MUX2 mux_inst_2 (
  .O(dout[0]),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(dff_q_0)
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(prom_inst_4_dout[1]),
  .I1(prom_inst_5_dout[1]),
  .S0(dff_q_1)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(prom_inst_6_dout[1]),
  .I1(prom_inst_7_dout[1]),
  .S0(dff_q_1)
);
MUX2 mux_inst_5 (
  .O(dout[1]),
  .I0(mux_o_3),
  .I1(mux_o_4),
  .S0(dff_q_0)
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(prom_inst_8_dout[2]),
  .I1(prom_inst_9_dout[2]),
  .S0(dff_q_1)
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(prom_inst_10_dout[2]),
  .I1(prom_inst_11_dout[2]),
  .S0(dff_q_1)
);
MUX2 mux_inst_8 (
  .O(dout[2]),
  .I0(mux_o_6),
  .I1(mux_o_7),
  .S0(dff_q_0)
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(prom_inst_12_dout[3]),
  .I1(prom_inst_13_dout[3]),
  .S0(dff_q_1)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(prom_inst_14_dout[3]),
  .I1(prom_inst_15_dout[3]),
  .S0(dff_q_1)
);
MUX2 mux_inst_11 (
  .O(dout[3]),
  .I0(mux_o_9),
  .I1(mux_o_10),
  .S0(dff_q_0)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(prom_inst_16_dout[4]),
  .I1(prom_inst_17_dout[4]),
  .S0(dff_q_1)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(prom_inst_18_dout[4]),
  .I1(prom_inst_19_dout[4]),
  .S0(dff_q_1)
);
MUX2 mux_inst_14 (
  .O(dout[4]),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(dff_q_0)
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(prom_inst_20_dout[5]),
  .I1(prom_inst_21_dout[5]),
  .S0(dff_q_1)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(prom_inst_22_dout[5]),
  .I1(prom_inst_23_dout[5]),
  .S0(dff_q_1)
);
MUX2 mux_inst_17 (
  .O(dout[5]),
  .I0(mux_o_15),
  .I1(mux_o_16),
  .S0(dff_q_0)
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(prom_inst_24_dout[6]),
  .I1(prom_inst_25_dout[6]),
  .S0(dff_q_1)
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(prom_inst_26_dout[6]),
  .I1(prom_inst_27_dout[6]),
  .S0(dff_q_1)
);
MUX2 mux_inst_20 (
  .O(dout[6]),
  .I0(mux_o_18),
  .I1(mux_o_19),
  .S0(dff_q_0)
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(prom_inst_28_dout[7]),
  .I1(prom_inst_29_dout[7]),
  .S0(dff_q_1)
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(prom_inst_30_dout[7]),
  .I1(prom_inst_31_dout[7]),
  .S0(dff_q_1)
);
MUX2 mux_inst_23 (
  .O(dout[7]),
  .I0(mux_o_21),
  .I1(mux_o_22),
  .S0(dff_q_0)
);
endmodule //Gowin_pROM
